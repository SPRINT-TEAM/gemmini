module cc_dir_ext( // @[:anonymous source@2.2]
  input  [9:0]   RW0_addr, // @[:anonymous source@3.4]
  input          RW0_clk, // @[:anonymous source@4.4]
  input  [127:0] RW0_wdata, // @[:anonymous source@5.4]
  output [127:0] RW0_rdata, // @[:anonymous source@6.4]
  input          RW0_en, // @[:anonymous source@7.4]
  input          RW0_wmode, // @[:anonymous source@8.4]
  input  [7:0]   RW0_wmask // @[:anonymous source@9.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_wdata; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_rdata; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@11.4]
  wire [9:0] mem_0_1_RW0_addr; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_wdata; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_rdata; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@12.4]
  wire [9:0] mem_0_2_RW0_addr; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_wdata; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_rdata; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@13.4]
  wire [9:0] mem_0_3_RW0_addr; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_wdata; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_rdata; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@14.4]
  wire [9:0] mem_0_4_RW0_addr; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_wdata; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_rdata; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@15.4]
  wire [9:0] mem_0_5_RW0_addr; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_wdata; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_rdata; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@16.4]
  wire [9:0] mem_0_6_RW0_addr; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_wdata; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_rdata; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@17.4]
  wire [9:0] mem_0_7_RW0_addr; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_wdata; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_rdata; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@18.4]
  wire [15:0] RW0_rdata_0_0; // @[:anonymous source@21.4]
  wire [15:0] RW0_rdata_0_1; // @[:anonymous source@28.4]
  wire [15:0] RW0_rdata_0_2; // @[:anonymous source@35.4]
  wire [15:0] RW0_rdata_0_3; // @[:anonymous source@42.4]
  wire [15:0] RW0_rdata_0_4; // @[:anonymous source@49.4]
  wire [15:0] RW0_rdata_0_5; // @[:anonymous source@56.4]
  wire [15:0] RW0_rdata_0_6; // @[:anonymous source@63.4]
  wire [15:0] RW0_rdata_0_7; // @[:anonymous source@70.4]
  wire [31:0] _GEN_0; // @[:anonymous source@75.4]
  wire [47:0] _GEN_1; // @[:anonymous source@75.4]
  wire [63:0] _GEN_2; // @[:anonymous source@75.4]
  wire [79:0] _GEN_3; // @[:anonymous source@75.4]
  wire [95:0] _GEN_4; // @[:anonymous source@75.4]
  wire [111:0] _GEN_5; // @[:anonymous source@75.4]
  wire [127:0] RW0_rdata_0; // @[:anonymous source@75.4]
  wire [31:0] _GEN_6; // @[:anonymous source@76.4]
  wire [47:0] _GEN_7; // @[:anonymous source@76.4]
  wire [63:0] _GEN_8; // @[:anonymous source@76.4]
  wire [79:0] _GEN_9; // @[:anonymous source@76.4]
  wire [95:0] _GEN_10; // @[:anonymous source@76.4]
  wire [111:0] _GEN_11; // @[:anonymous source@76.4]
  split_cc_dir_ext mem_0_0 ( // @[:anonymous source@11.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 ( // @[:anonymous source@12.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 ( // @[:anonymous source@13.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 ( // @[:anonymous source@14.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 ( // @[:anonymous source@15.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 ( // @[:anonymous source@16.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 ( // @[:anonymous source@17.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 ( // @[:anonymous source@18.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@21.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@28.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@35.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@42.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@49.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@56.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@63.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@70.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[:anonymous source@76.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@20.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@19.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[15:0]; // @[:anonymous source@22.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@25.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@24.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@23.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@27.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@26.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[31:16]; // @[:anonymous source@29.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@32.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@31.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@30.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@34.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@33.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[47:32]; // @[:anonymous source@36.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@39.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@38.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@37.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@41.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@40.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[63:48]; // @[:anonymous source@43.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@46.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@45.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@44.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@48.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@47.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[79:64]; // @[:anonymous source@50.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@53.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@52.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@51.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@55.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@54.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[95:80]; // @[:anonymous source@57.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@60.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@59.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@58.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@62.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@61.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[111:96]; // @[:anonymous source@64.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@67.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@66.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@65.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@69.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@68.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[127:112]; // @[:anonymous source@71.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@74.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@73.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@72.4]
endmodule
module cc_banks_0_ext( // @[:anonymous source@78.2]
  input  [12:0] RW0_addr, // @[:anonymous source@79.4]
  input         RW0_clk, // @[:anonymous source@80.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@81.4]
  output [63:0] RW0_rdata, // @[:anonymous source@82.4]
  input         RW0_en, // @[:anonymous source@83.4]
  input         RW0_wmode // @[:anonymous source@84.4]
);
  wire [12:0] mem_0_0_RW0_addr; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@86.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@89.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@93.4]
  split_cc_banks_0_ext mem_0_0 ( // @[:anonymous source@86.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@89.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@93.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@94.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@88.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@87.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@90.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@92.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@91.4]
endmodule
module data_arrays_0_ext( // @[:anonymous source@96.2]
  input  [7:0]   RW0_addr, // @[:anonymous source@97.4]
  input          RW0_clk, // @[:anonymous source@98.4]
  input  [255:0] RW0_wdata, // @[:anonymous source@99.4]
  output [255:0] RW0_rdata, // @[:anonymous source@100.4]
  input          RW0_en, // @[:anonymous source@101.4]
  input          RW0_wmode, // @[:anonymous source@102.4]
  input  [31:0]  RW0_wmask // @[:anonymous source@103.4]
);
  wire [7:0] mem_0_0_RW0_addr; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@105.4]
  wire [7:0] mem_0_0_RW0_wdata; // @[:anonymous source@105.4]
  wire [7:0] mem_0_0_RW0_rdata; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@105.4]
  wire [7:0] mem_0_1_RW0_addr; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@106.4]
  wire [7:0] mem_0_1_RW0_wdata; // @[:anonymous source@106.4]
  wire [7:0] mem_0_1_RW0_rdata; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@106.4]
  wire [7:0] mem_0_2_RW0_addr; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@107.4]
  wire [7:0] mem_0_2_RW0_wdata; // @[:anonymous source@107.4]
  wire [7:0] mem_0_2_RW0_rdata; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@107.4]
  wire [7:0] mem_0_3_RW0_addr; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@108.4]
  wire [7:0] mem_0_3_RW0_wdata; // @[:anonymous source@108.4]
  wire [7:0] mem_0_3_RW0_rdata; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@108.4]
  wire [7:0] mem_0_4_RW0_addr; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@109.4]
  wire [7:0] mem_0_4_RW0_wdata; // @[:anonymous source@109.4]
  wire [7:0] mem_0_4_RW0_rdata; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@109.4]
  wire [7:0] mem_0_5_RW0_addr; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@110.4]
  wire [7:0] mem_0_5_RW0_wdata; // @[:anonymous source@110.4]
  wire [7:0] mem_0_5_RW0_rdata; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@110.4]
  wire [7:0] mem_0_6_RW0_addr; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@111.4]
  wire [7:0] mem_0_6_RW0_wdata; // @[:anonymous source@111.4]
  wire [7:0] mem_0_6_RW0_rdata; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@111.4]
  wire [7:0] mem_0_7_RW0_addr; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@112.4]
  wire [7:0] mem_0_7_RW0_wdata; // @[:anonymous source@112.4]
  wire [7:0] mem_0_7_RW0_rdata; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@112.4]
  wire [7:0] mem_0_8_RW0_addr; // @[:anonymous source@113.4]
  wire  mem_0_8_RW0_clk; // @[:anonymous source@113.4]
  wire [7:0] mem_0_8_RW0_wdata; // @[:anonymous source@113.4]
  wire [7:0] mem_0_8_RW0_rdata; // @[:anonymous source@113.4]
  wire  mem_0_8_RW0_en; // @[:anonymous source@113.4]
  wire  mem_0_8_RW0_wmode; // @[:anonymous source@113.4]
  wire  mem_0_8_RW0_wmask; // @[:anonymous source@113.4]
  wire [7:0] mem_0_9_RW0_addr; // @[:anonymous source@114.4]
  wire  mem_0_9_RW0_clk; // @[:anonymous source@114.4]
  wire [7:0] mem_0_9_RW0_wdata; // @[:anonymous source@114.4]
  wire [7:0] mem_0_9_RW0_rdata; // @[:anonymous source@114.4]
  wire  mem_0_9_RW0_en; // @[:anonymous source@114.4]
  wire  mem_0_9_RW0_wmode; // @[:anonymous source@114.4]
  wire  mem_0_9_RW0_wmask; // @[:anonymous source@114.4]
  wire [7:0] mem_0_10_RW0_addr; // @[:anonymous source@115.4]
  wire  mem_0_10_RW0_clk; // @[:anonymous source@115.4]
  wire [7:0] mem_0_10_RW0_wdata; // @[:anonymous source@115.4]
  wire [7:0] mem_0_10_RW0_rdata; // @[:anonymous source@115.4]
  wire  mem_0_10_RW0_en; // @[:anonymous source@115.4]
  wire  mem_0_10_RW0_wmode; // @[:anonymous source@115.4]
  wire  mem_0_10_RW0_wmask; // @[:anonymous source@115.4]
  wire [7:0] mem_0_11_RW0_addr; // @[:anonymous source@116.4]
  wire  mem_0_11_RW0_clk; // @[:anonymous source@116.4]
  wire [7:0] mem_0_11_RW0_wdata; // @[:anonymous source@116.4]
  wire [7:0] mem_0_11_RW0_rdata; // @[:anonymous source@116.4]
  wire  mem_0_11_RW0_en; // @[:anonymous source@116.4]
  wire  mem_0_11_RW0_wmode; // @[:anonymous source@116.4]
  wire  mem_0_11_RW0_wmask; // @[:anonymous source@116.4]
  wire [7:0] mem_0_12_RW0_addr; // @[:anonymous source@117.4]
  wire  mem_0_12_RW0_clk; // @[:anonymous source@117.4]
  wire [7:0] mem_0_12_RW0_wdata; // @[:anonymous source@117.4]
  wire [7:0] mem_0_12_RW0_rdata; // @[:anonymous source@117.4]
  wire  mem_0_12_RW0_en; // @[:anonymous source@117.4]
  wire  mem_0_12_RW0_wmode; // @[:anonymous source@117.4]
  wire  mem_0_12_RW0_wmask; // @[:anonymous source@117.4]
  wire [7:0] mem_0_13_RW0_addr; // @[:anonymous source@118.4]
  wire  mem_0_13_RW0_clk; // @[:anonymous source@118.4]
  wire [7:0] mem_0_13_RW0_wdata; // @[:anonymous source@118.4]
  wire [7:0] mem_0_13_RW0_rdata; // @[:anonymous source@118.4]
  wire  mem_0_13_RW0_en; // @[:anonymous source@118.4]
  wire  mem_0_13_RW0_wmode; // @[:anonymous source@118.4]
  wire  mem_0_13_RW0_wmask; // @[:anonymous source@118.4]
  wire [7:0] mem_0_14_RW0_addr; // @[:anonymous source@119.4]
  wire  mem_0_14_RW0_clk; // @[:anonymous source@119.4]
  wire [7:0] mem_0_14_RW0_wdata; // @[:anonymous source@119.4]
  wire [7:0] mem_0_14_RW0_rdata; // @[:anonymous source@119.4]
  wire  mem_0_14_RW0_en; // @[:anonymous source@119.4]
  wire  mem_0_14_RW0_wmode; // @[:anonymous source@119.4]
  wire  mem_0_14_RW0_wmask; // @[:anonymous source@119.4]
  wire [7:0] mem_0_15_RW0_addr; // @[:anonymous source@120.4]
  wire  mem_0_15_RW0_clk; // @[:anonymous source@120.4]
  wire [7:0] mem_0_15_RW0_wdata; // @[:anonymous source@120.4]
  wire [7:0] mem_0_15_RW0_rdata; // @[:anonymous source@120.4]
  wire  mem_0_15_RW0_en; // @[:anonymous source@120.4]
  wire  mem_0_15_RW0_wmode; // @[:anonymous source@120.4]
  wire  mem_0_15_RW0_wmask; // @[:anonymous source@120.4]
  wire [7:0] mem_0_16_RW0_addr; // @[:anonymous source@121.4]
  wire  mem_0_16_RW0_clk; // @[:anonymous source@121.4]
  wire [7:0] mem_0_16_RW0_wdata; // @[:anonymous source@121.4]
  wire [7:0] mem_0_16_RW0_rdata; // @[:anonymous source@121.4]
  wire  mem_0_16_RW0_en; // @[:anonymous source@121.4]
  wire  mem_0_16_RW0_wmode; // @[:anonymous source@121.4]
  wire  mem_0_16_RW0_wmask; // @[:anonymous source@121.4]
  wire [7:0] mem_0_17_RW0_addr; // @[:anonymous source@122.4]
  wire  mem_0_17_RW0_clk; // @[:anonymous source@122.4]
  wire [7:0] mem_0_17_RW0_wdata; // @[:anonymous source@122.4]
  wire [7:0] mem_0_17_RW0_rdata; // @[:anonymous source@122.4]
  wire  mem_0_17_RW0_en; // @[:anonymous source@122.4]
  wire  mem_0_17_RW0_wmode; // @[:anonymous source@122.4]
  wire  mem_0_17_RW0_wmask; // @[:anonymous source@122.4]
  wire [7:0] mem_0_18_RW0_addr; // @[:anonymous source@123.4]
  wire  mem_0_18_RW0_clk; // @[:anonymous source@123.4]
  wire [7:0] mem_0_18_RW0_wdata; // @[:anonymous source@123.4]
  wire [7:0] mem_0_18_RW0_rdata; // @[:anonymous source@123.4]
  wire  mem_0_18_RW0_en; // @[:anonymous source@123.4]
  wire  mem_0_18_RW0_wmode; // @[:anonymous source@123.4]
  wire  mem_0_18_RW0_wmask; // @[:anonymous source@123.4]
  wire [7:0] mem_0_19_RW0_addr; // @[:anonymous source@124.4]
  wire  mem_0_19_RW0_clk; // @[:anonymous source@124.4]
  wire [7:0] mem_0_19_RW0_wdata; // @[:anonymous source@124.4]
  wire [7:0] mem_0_19_RW0_rdata; // @[:anonymous source@124.4]
  wire  mem_0_19_RW0_en; // @[:anonymous source@124.4]
  wire  mem_0_19_RW0_wmode; // @[:anonymous source@124.4]
  wire  mem_0_19_RW0_wmask; // @[:anonymous source@124.4]
  wire [7:0] mem_0_20_RW0_addr; // @[:anonymous source@125.4]
  wire  mem_0_20_RW0_clk; // @[:anonymous source@125.4]
  wire [7:0] mem_0_20_RW0_wdata; // @[:anonymous source@125.4]
  wire [7:0] mem_0_20_RW0_rdata; // @[:anonymous source@125.4]
  wire  mem_0_20_RW0_en; // @[:anonymous source@125.4]
  wire  mem_0_20_RW0_wmode; // @[:anonymous source@125.4]
  wire  mem_0_20_RW0_wmask; // @[:anonymous source@125.4]
  wire [7:0] mem_0_21_RW0_addr; // @[:anonymous source@126.4]
  wire  mem_0_21_RW0_clk; // @[:anonymous source@126.4]
  wire [7:0] mem_0_21_RW0_wdata; // @[:anonymous source@126.4]
  wire [7:0] mem_0_21_RW0_rdata; // @[:anonymous source@126.4]
  wire  mem_0_21_RW0_en; // @[:anonymous source@126.4]
  wire  mem_0_21_RW0_wmode; // @[:anonymous source@126.4]
  wire  mem_0_21_RW0_wmask; // @[:anonymous source@126.4]
  wire [7:0] mem_0_22_RW0_addr; // @[:anonymous source@127.4]
  wire  mem_0_22_RW0_clk; // @[:anonymous source@127.4]
  wire [7:0] mem_0_22_RW0_wdata; // @[:anonymous source@127.4]
  wire [7:0] mem_0_22_RW0_rdata; // @[:anonymous source@127.4]
  wire  mem_0_22_RW0_en; // @[:anonymous source@127.4]
  wire  mem_0_22_RW0_wmode; // @[:anonymous source@127.4]
  wire  mem_0_22_RW0_wmask; // @[:anonymous source@127.4]
  wire [7:0] mem_0_23_RW0_addr; // @[:anonymous source@128.4]
  wire  mem_0_23_RW0_clk; // @[:anonymous source@128.4]
  wire [7:0] mem_0_23_RW0_wdata; // @[:anonymous source@128.4]
  wire [7:0] mem_0_23_RW0_rdata; // @[:anonymous source@128.4]
  wire  mem_0_23_RW0_en; // @[:anonymous source@128.4]
  wire  mem_0_23_RW0_wmode; // @[:anonymous source@128.4]
  wire  mem_0_23_RW0_wmask; // @[:anonymous source@128.4]
  wire [7:0] mem_0_24_RW0_addr; // @[:anonymous source@129.4]
  wire  mem_0_24_RW0_clk; // @[:anonymous source@129.4]
  wire [7:0] mem_0_24_RW0_wdata; // @[:anonymous source@129.4]
  wire [7:0] mem_0_24_RW0_rdata; // @[:anonymous source@129.4]
  wire  mem_0_24_RW0_en; // @[:anonymous source@129.4]
  wire  mem_0_24_RW0_wmode; // @[:anonymous source@129.4]
  wire  mem_0_24_RW0_wmask; // @[:anonymous source@129.4]
  wire [7:0] mem_0_25_RW0_addr; // @[:anonymous source@130.4]
  wire  mem_0_25_RW0_clk; // @[:anonymous source@130.4]
  wire [7:0] mem_0_25_RW0_wdata; // @[:anonymous source@130.4]
  wire [7:0] mem_0_25_RW0_rdata; // @[:anonymous source@130.4]
  wire  mem_0_25_RW0_en; // @[:anonymous source@130.4]
  wire  mem_0_25_RW0_wmode; // @[:anonymous source@130.4]
  wire  mem_0_25_RW0_wmask; // @[:anonymous source@130.4]
  wire [7:0] mem_0_26_RW0_addr; // @[:anonymous source@131.4]
  wire  mem_0_26_RW0_clk; // @[:anonymous source@131.4]
  wire [7:0] mem_0_26_RW0_wdata; // @[:anonymous source@131.4]
  wire [7:0] mem_0_26_RW0_rdata; // @[:anonymous source@131.4]
  wire  mem_0_26_RW0_en; // @[:anonymous source@131.4]
  wire  mem_0_26_RW0_wmode; // @[:anonymous source@131.4]
  wire  mem_0_26_RW0_wmask; // @[:anonymous source@131.4]
  wire [7:0] mem_0_27_RW0_addr; // @[:anonymous source@132.4]
  wire  mem_0_27_RW0_clk; // @[:anonymous source@132.4]
  wire [7:0] mem_0_27_RW0_wdata; // @[:anonymous source@132.4]
  wire [7:0] mem_0_27_RW0_rdata; // @[:anonymous source@132.4]
  wire  mem_0_27_RW0_en; // @[:anonymous source@132.4]
  wire  mem_0_27_RW0_wmode; // @[:anonymous source@132.4]
  wire  mem_0_27_RW0_wmask; // @[:anonymous source@132.4]
  wire [7:0] mem_0_28_RW0_addr; // @[:anonymous source@133.4]
  wire  mem_0_28_RW0_clk; // @[:anonymous source@133.4]
  wire [7:0] mem_0_28_RW0_wdata; // @[:anonymous source@133.4]
  wire [7:0] mem_0_28_RW0_rdata; // @[:anonymous source@133.4]
  wire  mem_0_28_RW0_en; // @[:anonymous source@133.4]
  wire  mem_0_28_RW0_wmode; // @[:anonymous source@133.4]
  wire  mem_0_28_RW0_wmask; // @[:anonymous source@133.4]
  wire [7:0] mem_0_29_RW0_addr; // @[:anonymous source@134.4]
  wire  mem_0_29_RW0_clk; // @[:anonymous source@134.4]
  wire [7:0] mem_0_29_RW0_wdata; // @[:anonymous source@134.4]
  wire [7:0] mem_0_29_RW0_rdata; // @[:anonymous source@134.4]
  wire  mem_0_29_RW0_en; // @[:anonymous source@134.4]
  wire  mem_0_29_RW0_wmode; // @[:anonymous source@134.4]
  wire  mem_0_29_RW0_wmask; // @[:anonymous source@134.4]
  wire [7:0] mem_0_30_RW0_addr; // @[:anonymous source@135.4]
  wire  mem_0_30_RW0_clk; // @[:anonymous source@135.4]
  wire [7:0] mem_0_30_RW0_wdata; // @[:anonymous source@135.4]
  wire [7:0] mem_0_30_RW0_rdata; // @[:anonymous source@135.4]
  wire  mem_0_30_RW0_en; // @[:anonymous source@135.4]
  wire  mem_0_30_RW0_wmode; // @[:anonymous source@135.4]
  wire  mem_0_30_RW0_wmask; // @[:anonymous source@135.4]
  wire [7:0] mem_0_31_RW0_addr; // @[:anonymous source@136.4]
  wire  mem_0_31_RW0_clk; // @[:anonymous source@136.4]
  wire [7:0] mem_0_31_RW0_wdata; // @[:anonymous source@136.4]
  wire [7:0] mem_0_31_RW0_rdata; // @[:anonymous source@136.4]
  wire  mem_0_31_RW0_en; // @[:anonymous source@136.4]
  wire  mem_0_31_RW0_wmode; // @[:anonymous source@136.4]
  wire  mem_0_31_RW0_wmask; // @[:anonymous source@136.4]
  wire [7:0] RW0_rdata_0_0; // @[:anonymous source@139.4]
  wire [7:0] RW0_rdata_0_1; // @[:anonymous source@146.4]
  wire [7:0] RW0_rdata_0_2; // @[:anonymous source@153.4]
  wire [7:0] RW0_rdata_0_3; // @[:anonymous source@160.4]
  wire [7:0] RW0_rdata_0_4; // @[:anonymous source@167.4]
  wire [7:0] RW0_rdata_0_5; // @[:anonymous source@174.4]
  wire [7:0] RW0_rdata_0_6; // @[:anonymous source@181.4]
  wire [7:0] RW0_rdata_0_7; // @[:anonymous source@188.4]
  wire [7:0] RW0_rdata_0_8; // @[:anonymous source@195.4]
  wire [7:0] RW0_rdata_0_9; // @[:anonymous source@202.4]
  wire [7:0] RW0_rdata_0_10; // @[:anonymous source@209.4]
  wire [7:0] RW0_rdata_0_11; // @[:anonymous source@216.4]
  wire [7:0] RW0_rdata_0_12; // @[:anonymous source@223.4]
  wire [7:0] RW0_rdata_0_13; // @[:anonymous source@230.4]
  wire [7:0] RW0_rdata_0_14; // @[:anonymous source@237.4]
  wire [7:0] RW0_rdata_0_15; // @[:anonymous source@244.4]
  wire [7:0] RW0_rdata_0_16; // @[:anonymous source@251.4]
  wire [7:0] RW0_rdata_0_17; // @[:anonymous source@258.4]
  wire [7:0] RW0_rdata_0_18; // @[:anonymous source@265.4]
  wire [7:0] RW0_rdata_0_19; // @[:anonymous source@272.4]
  wire [7:0] RW0_rdata_0_20; // @[:anonymous source@279.4]
  wire [7:0] RW0_rdata_0_21; // @[:anonymous source@286.4]
  wire [7:0] RW0_rdata_0_22; // @[:anonymous source@293.4]
  wire [7:0] RW0_rdata_0_23; // @[:anonymous source@300.4]
  wire [7:0] RW0_rdata_0_24; // @[:anonymous source@307.4]
  wire [7:0] RW0_rdata_0_25; // @[:anonymous source@314.4]
  wire [7:0] RW0_rdata_0_26; // @[:anonymous source@321.4]
  wire [7:0] RW0_rdata_0_27; // @[:anonymous source@328.4]
  wire [7:0] RW0_rdata_0_28; // @[:anonymous source@335.4]
  wire [7:0] RW0_rdata_0_29; // @[:anonymous source@342.4]
  wire [7:0] RW0_rdata_0_30; // @[:anonymous source@349.4]
  wire [7:0] RW0_rdata_0_31; // @[:anonymous source@356.4]
  wire [15:0] _GEN_0; // @[:anonymous source@361.4]
  wire [23:0] _GEN_1; // @[:anonymous source@361.4]
  wire [31:0] _GEN_2; // @[:anonymous source@361.4]
  wire [39:0] _GEN_3; // @[:anonymous source@361.4]
  wire [47:0] _GEN_4; // @[:anonymous source@361.4]
  wire [55:0] _GEN_5; // @[:anonymous source@361.4]
  wire [63:0] _GEN_6; // @[:anonymous source@361.4]
  wire [71:0] _GEN_7; // @[:anonymous source@361.4]
  wire [79:0] _GEN_8; // @[:anonymous source@361.4]
  wire [87:0] _GEN_9; // @[:anonymous source@361.4]
  wire [95:0] _GEN_10; // @[:anonymous source@361.4]
  wire [103:0] _GEN_11; // @[:anonymous source@361.4]
  wire [111:0] _GEN_12; // @[:anonymous source@361.4]
  wire [119:0] _GEN_13; // @[:anonymous source@361.4]
  wire [127:0] _GEN_14; // @[:anonymous source@361.4]
  wire [135:0] _GEN_15; // @[:anonymous source@361.4]
  wire [143:0] _GEN_16; // @[:anonymous source@361.4]
  wire [151:0] _GEN_17; // @[:anonymous source@361.4]
  wire [159:0] _GEN_18; // @[:anonymous source@361.4]
  wire [167:0] _GEN_19; // @[:anonymous source@361.4]
  wire [175:0] _GEN_20; // @[:anonymous source@361.4]
  wire [183:0] _GEN_21; // @[:anonymous source@361.4]
  wire [191:0] _GEN_22; // @[:anonymous source@361.4]
  wire [199:0] _GEN_23; // @[:anonymous source@361.4]
  wire [207:0] _GEN_24; // @[:anonymous source@361.4]
  wire [215:0] _GEN_25; // @[:anonymous source@361.4]
  wire [223:0] _GEN_26; // @[:anonymous source@361.4]
  wire [231:0] _GEN_27; // @[:anonymous source@361.4]
  wire [239:0] _GEN_28; // @[:anonymous source@361.4]
  wire [247:0] _GEN_29; // @[:anonymous source@361.4]
  wire [255:0] RW0_rdata_0; // @[:anonymous source@361.4]
  wire [15:0] _GEN_30; // @[:anonymous source@362.4]
  wire [23:0] _GEN_31; // @[:anonymous source@362.4]
  wire [31:0] _GEN_32; // @[:anonymous source@362.4]
  wire [39:0] _GEN_33; // @[:anonymous source@362.4]
  wire [47:0] _GEN_34; // @[:anonymous source@362.4]
  wire [55:0] _GEN_35; // @[:anonymous source@362.4]
  wire [63:0] _GEN_36; // @[:anonymous source@362.4]
  wire [71:0] _GEN_37; // @[:anonymous source@362.4]
  wire [79:0] _GEN_38; // @[:anonymous source@362.4]
  wire [87:0] _GEN_39; // @[:anonymous source@362.4]
  wire [95:0] _GEN_40; // @[:anonymous source@362.4]
  wire [103:0] _GEN_41; // @[:anonymous source@362.4]
  wire [111:0] _GEN_42; // @[:anonymous source@362.4]
  wire [119:0] _GEN_43; // @[:anonymous source@362.4]
  wire [127:0] _GEN_44; // @[:anonymous source@362.4]
  wire [135:0] _GEN_45; // @[:anonymous source@362.4]
  wire [143:0] _GEN_46; // @[:anonymous source@362.4]
  wire [151:0] _GEN_47; // @[:anonymous source@362.4]
  wire [159:0] _GEN_48; // @[:anonymous source@362.4]
  wire [167:0] _GEN_49; // @[:anonymous source@362.4]
  wire [175:0] _GEN_50; // @[:anonymous source@362.4]
  wire [183:0] _GEN_51; // @[:anonymous source@362.4]
  wire [191:0] _GEN_52; // @[:anonymous source@362.4]
  wire [199:0] _GEN_53; // @[:anonymous source@362.4]
  wire [207:0] _GEN_54; // @[:anonymous source@362.4]
  wire [215:0] _GEN_55; // @[:anonymous source@362.4]
  wire [223:0] _GEN_56; // @[:anonymous source@362.4]
  wire [231:0] _GEN_57; // @[:anonymous source@362.4]
  wire [239:0] _GEN_58; // @[:anonymous source@362.4]
  wire [247:0] _GEN_59; // @[:anonymous source@362.4]
  split_data_arrays_0_ext mem_0_0 ( // @[:anonymous source@105.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_1 ( // @[:anonymous source@106.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_2 ( // @[:anonymous source@107.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_3 ( // @[:anonymous source@108.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_4 ( // @[:anonymous source@109.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_5 ( // @[:anonymous source@110.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_6 ( // @[:anonymous source@111.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_7 ( // @[:anonymous source@112.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_8 ( // @[:anonymous source@113.4]
    .RW0_addr(mem_0_8_RW0_addr),
    .RW0_clk(mem_0_8_RW0_clk),
    .RW0_wdata(mem_0_8_RW0_wdata),
    .RW0_rdata(mem_0_8_RW0_rdata),
    .RW0_en(mem_0_8_RW0_en),
    .RW0_wmode(mem_0_8_RW0_wmode),
    .RW0_wmask(mem_0_8_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_9 ( // @[:anonymous source@114.4]
    .RW0_addr(mem_0_9_RW0_addr),
    .RW0_clk(mem_0_9_RW0_clk),
    .RW0_wdata(mem_0_9_RW0_wdata),
    .RW0_rdata(mem_0_9_RW0_rdata),
    .RW0_en(mem_0_9_RW0_en),
    .RW0_wmode(mem_0_9_RW0_wmode),
    .RW0_wmask(mem_0_9_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_10 ( // @[:anonymous source@115.4]
    .RW0_addr(mem_0_10_RW0_addr),
    .RW0_clk(mem_0_10_RW0_clk),
    .RW0_wdata(mem_0_10_RW0_wdata),
    .RW0_rdata(mem_0_10_RW0_rdata),
    .RW0_en(mem_0_10_RW0_en),
    .RW0_wmode(mem_0_10_RW0_wmode),
    .RW0_wmask(mem_0_10_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_11 ( // @[:anonymous source@116.4]
    .RW0_addr(mem_0_11_RW0_addr),
    .RW0_clk(mem_0_11_RW0_clk),
    .RW0_wdata(mem_0_11_RW0_wdata),
    .RW0_rdata(mem_0_11_RW0_rdata),
    .RW0_en(mem_0_11_RW0_en),
    .RW0_wmode(mem_0_11_RW0_wmode),
    .RW0_wmask(mem_0_11_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_12 ( // @[:anonymous source@117.4]
    .RW0_addr(mem_0_12_RW0_addr),
    .RW0_clk(mem_0_12_RW0_clk),
    .RW0_wdata(mem_0_12_RW0_wdata),
    .RW0_rdata(mem_0_12_RW0_rdata),
    .RW0_en(mem_0_12_RW0_en),
    .RW0_wmode(mem_0_12_RW0_wmode),
    .RW0_wmask(mem_0_12_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_13 ( // @[:anonymous source@118.4]
    .RW0_addr(mem_0_13_RW0_addr),
    .RW0_clk(mem_0_13_RW0_clk),
    .RW0_wdata(mem_0_13_RW0_wdata),
    .RW0_rdata(mem_0_13_RW0_rdata),
    .RW0_en(mem_0_13_RW0_en),
    .RW0_wmode(mem_0_13_RW0_wmode),
    .RW0_wmask(mem_0_13_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_14 ( // @[:anonymous source@119.4]
    .RW0_addr(mem_0_14_RW0_addr),
    .RW0_clk(mem_0_14_RW0_clk),
    .RW0_wdata(mem_0_14_RW0_wdata),
    .RW0_rdata(mem_0_14_RW0_rdata),
    .RW0_en(mem_0_14_RW0_en),
    .RW0_wmode(mem_0_14_RW0_wmode),
    .RW0_wmask(mem_0_14_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_15 ( // @[:anonymous source@120.4]
    .RW0_addr(mem_0_15_RW0_addr),
    .RW0_clk(mem_0_15_RW0_clk),
    .RW0_wdata(mem_0_15_RW0_wdata),
    .RW0_rdata(mem_0_15_RW0_rdata),
    .RW0_en(mem_0_15_RW0_en),
    .RW0_wmode(mem_0_15_RW0_wmode),
    .RW0_wmask(mem_0_15_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_16 ( // @[:anonymous source@121.4]
    .RW0_addr(mem_0_16_RW0_addr),
    .RW0_clk(mem_0_16_RW0_clk),
    .RW0_wdata(mem_0_16_RW0_wdata),
    .RW0_rdata(mem_0_16_RW0_rdata),
    .RW0_en(mem_0_16_RW0_en),
    .RW0_wmode(mem_0_16_RW0_wmode),
    .RW0_wmask(mem_0_16_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_17 ( // @[:anonymous source@122.4]
    .RW0_addr(mem_0_17_RW0_addr),
    .RW0_clk(mem_0_17_RW0_clk),
    .RW0_wdata(mem_0_17_RW0_wdata),
    .RW0_rdata(mem_0_17_RW0_rdata),
    .RW0_en(mem_0_17_RW0_en),
    .RW0_wmode(mem_0_17_RW0_wmode),
    .RW0_wmask(mem_0_17_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_18 ( // @[:anonymous source@123.4]
    .RW0_addr(mem_0_18_RW0_addr),
    .RW0_clk(mem_0_18_RW0_clk),
    .RW0_wdata(mem_0_18_RW0_wdata),
    .RW0_rdata(mem_0_18_RW0_rdata),
    .RW0_en(mem_0_18_RW0_en),
    .RW0_wmode(mem_0_18_RW0_wmode),
    .RW0_wmask(mem_0_18_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_19 ( // @[:anonymous source@124.4]
    .RW0_addr(mem_0_19_RW0_addr),
    .RW0_clk(mem_0_19_RW0_clk),
    .RW0_wdata(mem_0_19_RW0_wdata),
    .RW0_rdata(mem_0_19_RW0_rdata),
    .RW0_en(mem_0_19_RW0_en),
    .RW0_wmode(mem_0_19_RW0_wmode),
    .RW0_wmask(mem_0_19_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_20 ( // @[:anonymous source@125.4]
    .RW0_addr(mem_0_20_RW0_addr),
    .RW0_clk(mem_0_20_RW0_clk),
    .RW0_wdata(mem_0_20_RW0_wdata),
    .RW0_rdata(mem_0_20_RW0_rdata),
    .RW0_en(mem_0_20_RW0_en),
    .RW0_wmode(mem_0_20_RW0_wmode),
    .RW0_wmask(mem_0_20_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_21 ( // @[:anonymous source@126.4]
    .RW0_addr(mem_0_21_RW0_addr),
    .RW0_clk(mem_0_21_RW0_clk),
    .RW0_wdata(mem_0_21_RW0_wdata),
    .RW0_rdata(mem_0_21_RW0_rdata),
    .RW0_en(mem_0_21_RW0_en),
    .RW0_wmode(mem_0_21_RW0_wmode),
    .RW0_wmask(mem_0_21_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_22 ( // @[:anonymous source@127.4]
    .RW0_addr(mem_0_22_RW0_addr),
    .RW0_clk(mem_0_22_RW0_clk),
    .RW0_wdata(mem_0_22_RW0_wdata),
    .RW0_rdata(mem_0_22_RW0_rdata),
    .RW0_en(mem_0_22_RW0_en),
    .RW0_wmode(mem_0_22_RW0_wmode),
    .RW0_wmask(mem_0_22_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_23 ( // @[:anonymous source@128.4]
    .RW0_addr(mem_0_23_RW0_addr),
    .RW0_clk(mem_0_23_RW0_clk),
    .RW0_wdata(mem_0_23_RW0_wdata),
    .RW0_rdata(mem_0_23_RW0_rdata),
    .RW0_en(mem_0_23_RW0_en),
    .RW0_wmode(mem_0_23_RW0_wmode),
    .RW0_wmask(mem_0_23_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_24 ( // @[:anonymous source@129.4]
    .RW0_addr(mem_0_24_RW0_addr),
    .RW0_clk(mem_0_24_RW0_clk),
    .RW0_wdata(mem_0_24_RW0_wdata),
    .RW0_rdata(mem_0_24_RW0_rdata),
    .RW0_en(mem_0_24_RW0_en),
    .RW0_wmode(mem_0_24_RW0_wmode),
    .RW0_wmask(mem_0_24_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_25 ( // @[:anonymous source@130.4]
    .RW0_addr(mem_0_25_RW0_addr),
    .RW0_clk(mem_0_25_RW0_clk),
    .RW0_wdata(mem_0_25_RW0_wdata),
    .RW0_rdata(mem_0_25_RW0_rdata),
    .RW0_en(mem_0_25_RW0_en),
    .RW0_wmode(mem_0_25_RW0_wmode),
    .RW0_wmask(mem_0_25_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_26 ( // @[:anonymous source@131.4]
    .RW0_addr(mem_0_26_RW0_addr),
    .RW0_clk(mem_0_26_RW0_clk),
    .RW0_wdata(mem_0_26_RW0_wdata),
    .RW0_rdata(mem_0_26_RW0_rdata),
    .RW0_en(mem_0_26_RW0_en),
    .RW0_wmode(mem_0_26_RW0_wmode),
    .RW0_wmask(mem_0_26_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_27 ( // @[:anonymous source@132.4]
    .RW0_addr(mem_0_27_RW0_addr),
    .RW0_clk(mem_0_27_RW0_clk),
    .RW0_wdata(mem_0_27_RW0_wdata),
    .RW0_rdata(mem_0_27_RW0_rdata),
    .RW0_en(mem_0_27_RW0_en),
    .RW0_wmode(mem_0_27_RW0_wmode),
    .RW0_wmask(mem_0_27_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_28 ( // @[:anonymous source@133.4]
    .RW0_addr(mem_0_28_RW0_addr),
    .RW0_clk(mem_0_28_RW0_clk),
    .RW0_wdata(mem_0_28_RW0_wdata),
    .RW0_rdata(mem_0_28_RW0_rdata),
    .RW0_en(mem_0_28_RW0_en),
    .RW0_wmode(mem_0_28_RW0_wmode),
    .RW0_wmask(mem_0_28_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_29 ( // @[:anonymous source@134.4]
    .RW0_addr(mem_0_29_RW0_addr),
    .RW0_clk(mem_0_29_RW0_clk),
    .RW0_wdata(mem_0_29_RW0_wdata),
    .RW0_rdata(mem_0_29_RW0_rdata),
    .RW0_en(mem_0_29_RW0_en),
    .RW0_wmode(mem_0_29_RW0_wmode),
    .RW0_wmask(mem_0_29_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_30 ( // @[:anonymous source@135.4]
    .RW0_addr(mem_0_30_RW0_addr),
    .RW0_clk(mem_0_30_RW0_clk),
    .RW0_wdata(mem_0_30_RW0_wdata),
    .RW0_rdata(mem_0_30_RW0_rdata),
    .RW0_en(mem_0_30_RW0_en),
    .RW0_wmode(mem_0_30_RW0_wmode),
    .RW0_wmask(mem_0_30_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_31 ( // @[:anonymous source@136.4]
    .RW0_addr(mem_0_31_RW0_addr),
    .RW0_clk(mem_0_31_RW0_clk),
    .RW0_wdata(mem_0_31_RW0_wdata),
    .RW0_rdata(mem_0_31_RW0_rdata),
    .RW0_en(mem_0_31_RW0_en),
    .RW0_wmode(mem_0_31_RW0_wmode),
    .RW0_wmask(mem_0_31_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@139.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@146.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@153.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@160.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@167.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@174.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@181.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@188.4]
  assign RW0_rdata_0_8 = mem_0_8_RW0_rdata; // @[:anonymous source@195.4]
  assign RW0_rdata_0_9 = mem_0_9_RW0_rdata; // @[:anonymous source@202.4]
  assign RW0_rdata_0_10 = mem_0_10_RW0_rdata; // @[:anonymous source@209.4]
  assign RW0_rdata_0_11 = mem_0_11_RW0_rdata; // @[:anonymous source@216.4]
  assign RW0_rdata_0_12 = mem_0_12_RW0_rdata; // @[:anonymous source@223.4]
  assign RW0_rdata_0_13 = mem_0_13_RW0_rdata; // @[:anonymous source@230.4]
  assign RW0_rdata_0_14 = mem_0_14_RW0_rdata; // @[:anonymous source@237.4]
  assign RW0_rdata_0_15 = mem_0_15_RW0_rdata; // @[:anonymous source@244.4]
  assign RW0_rdata_0_16 = mem_0_16_RW0_rdata; // @[:anonymous source@251.4]
  assign RW0_rdata_0_17 = mem_0_17_RW0_rdata; // @[:anonymous source@258.4]
  assign RW0_rdata_0_18 = mem_0_18_RW0_rdata; // @[:anonymous source@265.4]
  assign RW0_rdata_0_19 = mem_0_19_RW0_rdata; // @[:anonymous source@272.4]
  assign RW0_rdata_0_20 = mem_0_20_RW0_rdata; // @[:anonymous source@279.4]
  assign RW0_rdata_0_21 = mem_0_21_RW0_rdata; // @[:anonymous source@286.4]
  assign RW0_rdata_0_22 = mem_0_22_RW0_rdata; // @[:anonymous source@293.4]
  assign RW0_rdata_0_23 = mem_0_23_RW0_rdata; // @[:anonymous source@300.4]
  assign RW0_rdata_0_24 = mem_0_24_RW0_rdata; // @[:anonymous source@307.4]
  assign RW0_rdata_0_25 = mem_0_25_RW0_rdata; // @[:anonymous source@314.4]
  assign RW0_rdata_0_26 = mem_0_26_RW0_rdata; // @[:anonymous source@321.4]
  assign RW0_rdata_0_27 = mem_0_27_RW0_rdata; // @[:anonymous source@328.4]
  assign RW0_rdata_0_28 = mem_0_28_RW0_rdata; // @[:anonymous source@335.4]
  assign RW0_rdata_0_29 = mem_0_29_RW0_rdata; // @[:anonymous source@342.4]
  assign RW0_rdata_0_30 = mem_0_30_RW0_rdata; // @[:anonymous source@349.4]
  assign RW0_rdata_0_31 = mem_0_31_RW0_rdata; // @[:anonymous source@356.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_6 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_7 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_8 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@361.4]
  assign _GEN_9 = {RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_10 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_11 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_12 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_13 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_14 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_15 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_16 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_17 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@361.4]
  assign _GEN_18 = {RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_19 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_20 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_21 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_22 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_23 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_24 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_25 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_26 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@361.4]
  assign _GEN_27 = {RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@361.4]
  assign _GEN_28 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@361.4]
  assign _GEN_29 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@361.4]
  assign RW0_rdata_0 = {RW0_rdata_0_31,RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@361.4]
  assign _GEN_30 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_31 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_32 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_33 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_34 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_35 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_36 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_37 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_38 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@362.4]
  assign _GEN_39 = {RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_40 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_41 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_42 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_43 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_44 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_45 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_46 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_47 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[:anonymous source@362.4]
  assign _GEN_48 = {RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_49 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_50 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_51 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_52 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_53 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_54 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_55 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_56 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[:anonymous source@362.4]
  assign _GEN_57 = {RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@362.4]
  assign _GEN_58 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@362.4]
  assign _GEN_59 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[:anonymous source@362.4]
  assign RW0_rdata = {RW0_rdata_0_31,_GEN_29}; // @[:anonymous source@362.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@138.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@137.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0]; // @[:anonymous source@140.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@143.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@142.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@141.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@145.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@144.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8]; // @[:anonymous source@147.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@150.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@149.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@148.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@152.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@151.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16]; // @[:anonymous source@154.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@157.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@156.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@155.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@159.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@158.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24]; // @[:anonymous source@161.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@164.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@163.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@162.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@166.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@165.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32]; // @[:anonymous source@168.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@171.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@170.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@169.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@173.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@172.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40]; // @[:anonymous source@175.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@178.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@177.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@176.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@180.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@179.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48]; // @[:anonymous source@182.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@185.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@184.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@183.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@187.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@186.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56]; // @[:anonymous source@189.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@192.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@191.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@190.4]
  assign mem_0_8_RW0_addr = RW0_addr; // @[:anonymous source@194.4]
  assign mem_0_8_RW0_clk = RW0_clk; // @[:anonymous source@193.4]
  assign mem_0_8_RW0_wdata = RW0_wdata[71:64]; // @[:anonymous source@196.4]
  assign mem_0_8_RW0_en = RW0_en; // @[:anonymous source@199.4]
  assign mem_0_8_RW0_wmode = RW0_wmode; // @[:anonymous source@198.4]
  assign mem_0_8_RW0_wmask = RW0_wmask[8]; // @[:anonymous source@197.4]
  assign mem_0_9_RW0_addr = RW0_addr; // @[:anonymous source@201.4]
  assign mem_0_9_RW0_clk = RW0_clk; // @[:anonymous source@200.4]
  assign mem_0_9_RW0_wdata = RW0_wdata[79:72]; // @[:anonymous source@203.4]
  assign mem_0_9_RW0_en = RW0_en; // @[:anonymous source@206.4]
  assign mem_0_9_RW0_wmode = RW0_wmode; // @[:anonymous source@205.4]
  assign mem_0_9_RW0_wmask = RW0_wmask[9]; // @[:anonymous source@204.4]
  assign mem_0_10_RW0_addr = RW0_addr; // @[:anonymous source@208.4]
  assign mem_0_10_RW0_clk = RW0_clk; // @[:anonymous source@207.4]
  assign mem_0_10_RW0_wdata = RW0_wdata[87:80]; // @[:anonymous source@210.4]
  assign mem_0_10_RW0_en = RW0_en; // @[:anonymous source@213.4]
  assign mem_0_10_RW0_wmode = RW0_wmode; // @[:anonymous source@212.4]
  assign mem_0_10_RW0_wmask = RW0_wmask[10]; // @[:anonymous source@211.4]
  assign mem_0_11_RW0_addr = RW0_addr; // @[:anonymous source@215.4]
  assign mem_0_11_RW0_clk = RW0_clk; // @[:anonymous source@214.4]
  assign mem_0_11_RW0_wdata = RW0_wdata[95:88]; // @[:anonymous source@217.4]
  assign mem_0_11_RW0_en = RW0_en; // @[:anonymous source@220.4]
  assign mem_0_11_RW0_wmode = RW0_wmode; // @[:anonymous source@219.4]
  assign mem_0_11_RW0_wmask = RW0_wmask[11]; // @[:anonymous source@218.4]
  assign mem_0_12_RW0_addr = RW0_addr; // @[:anonymous source@222.4]
  assign mem_0_12_RW0_clk = RW0_clk; // @[:anonymous source@221.4]
  assign mem_0_12_RW0_wdata = RW0_wdata[103:96]; // @[:anonymous source@224.4]
  assign mem_0_12_RW0_en = RW0_en; // @[:anonymous source@227.4]
  assign mem_0_12_RW0_wmode = RW0_wmode; // @[:anonymous source@226.4]
  assign mem_0_12_RW0_wmask = RW0_wmask[12]; // @[:anonymous source@225.4]
  assign mem_0_13_RW0_addr = RW0_addr; // @[:anonymous source@229.4]
  assign mem_0_13_RW0_clk = RW0_clk; // @[:anonymous source@228.4]
  assign mem_0_13_RW0_wdata = RW0_wdata[111:104]; // @[:anonymous source@231.4]
  assign mem_0_13_RW0_en = RW0_en; // @[:anonymous source@234.4]
  assign mem_0_13_RW0_wmode = RW0_wmode; // @[:anonymous source@233.4]
  assign mem_0_13_RW0_wmask = RW0_wmask[13]; // @[:anonymous source@232.4]
  assign mem_0_14_RW0_addr = RW0_addr; // @[:anonymous source@236.4]
  assign mem_0_14_RW0_clk = RW0_clk; // @[:anonymous source@235.4]
  assign mem_0_14_RW0_wdata = RW0_wdata[119:112]; // @[:anonymous source@238.4]
  assign mem_0_14_RW0_en = RW0_en; // @[:anonymous source@241.4]
  assign mem_0_14_RW0_wmode = RW0_wmode; // @[:anonymous source@240.4]
  assign mem_0_14_RW0_wmask = RW0_wmask[14]; // @[:anonymous source@239.4]
  assign mem_0_15_RW0_addr = RW0_addr; // @[:anonymous source@243.4]
  assign mem_0_15_RW0_clk = RW0_clk; // @[:anonymous source@242.4]
  assign mem_0_15_RW0_wdata = RW0_wdata[127:120]; // @[:anonymous source@245.4]
  assign mem_0_15_RW0_en = RW0_en; // @[:anonymous source@248.4]
  assign mem_0_15_RW0_wmode = RW0_wmode; // @[:anonymous source@247.4]
  assign mem_0_15_RW0_wmask = RW0_wmask[15]; // @[:anonymous source@246.4]
  assign mem_0_16_RW0_addr = RW0_addr; // @[:anonymous source@250.4]
  assign mem_0_16_RW0_clk = RW0_clk; // @[:anonymous source@249.4]
  assign mem_0_16_RW0_wdata = RW0_wdata[135:128]; // @[:anonymous source@252.4]
  assign mem_0_16_RW0_en = RW0_en; // @[:anonymous source@255.4]
  assign mem_0_16_RW0_wmode = RW0_wmode; // @[:anonymous source@254.4]
  assign mem_0_16_RW0_wmask = RW0_wmask[16]; // @[:anonymous source@253.4]
  assign mem_0_17_RW0_addr = RW0_addr; // @[:anonymous source@257.4]
  assign mem_0_17_RW0_clk = RW0_clk; // @[:anonymous source@256.4]
  assign mem_0_17_RW0_wdata = RW0_wdata[143:136]; // @[:anonymous source@259.4]
  assign mem_0_17_RW0_en = RW0_en; // @[:anonymous source@262.4]
  assign mem_0_17_RW0_wmode = RW0_wmode; // @[:anonymous source@261.4]
  assign mem_0_17_RW0_wmask = RW0_wmask[17]; // @[:anonymous source@260.4]
  assign mem_0_18_RW0_addr = RW0_addr; // @[:anonymous source@264.4]
  assign mem_0_18_RW0_clk = RW0_clk; // @[:anonymous source@263.4]
  assign mem_0_18_RW0_wdata = RW0_wdata[151:144]; // @[:anonymous source@266.4]
  assign mem_0_18_RW0_en = RW0_en; // @[:anonymous source@269.4]
  assign mem_0_18_RW0_wmode = RW0_wmode; // @[:anonymous source@268.4]
  assign mem_0_18_RW0_wmask = RW0_wmask[18]; // @[:anonymous source@267.4]
  assign mem_0_19_RW0_addr = RW0_addr; // @[:anonymous source@271.4]
  assign mem_0_19_RW0_clk = RW0_clk; // @[:anonymous source@270.4]
  assign mem_0_19_RW0_wdata = RW0_wdata[159:152]; // @[:anonymous source@273.4]
  assign mem_0_19_RW0_en = RW0_en; // @[:anonymous source@276.4]
  assign mem_0_19_RW0_wmode = RW0_wmode; // @[:anonymous source@275.4]
  assign mem_0_19_RW0_wmask = RW0_wmask[19]; // @[:anonymous source@274.4]
  assign mem_0_20_RW0_addr = RW0_addr; // @[:anonymous source@278.4]
  assign mem_0_20_RW0_clk = RW0_clk; // @[:anonymous source@277.4]
  assign mem_0_20_RW0_wdata = RW0_wdata[167:160]; // @[:anonymous source@280.4]
  assign mem_0_20_RW0_en = RW0_en; // @[:anonymous source@283.4]
  assign mem_0_20_RW0_wmode = RW0_wmode; // @[:anonymous source@282.4]
  assign mem_0_20_RW0_wmask = RW0_wmask[20]; // @[:anonymous source@281.4]
  assign mem_0_21_RW0_addr = RW0_addr; // @[:anonymous source@285.4]
  assign mem_0_21_RW0_clk = RW0_clk; // @[:anonymous source@284.4]
  assign mem_0_21_RW0_wdata = RW0_wdata[175:168]; // @[:anonymous source@287.4]
  assign mem_0_21_RW0_en = RW0_en; // @[:anonymous source@290.4]
  assign mem_0_21_RW0_wmode = RW0_wmode; // @[:anonymous source@289.4]
  assign mem_0_21_RW0_wmask = RW0_wmask[21]; // @[:anonymous source@288.4]
  assign mem_0_22_RW0_addr = RW0_addr; // @[:anonymous source@292.4]
  assign mem_0_22_RW0_clk = RW0_clk; // @[:anonymous source@291.4]
  assign mem_0_22_RW0_wdata = RW0_wdata[183:176]; // @[:anonymous source@294.4]
  assign mem_0_22_RW0_en = RW0_en; // @[:anonymous source@297.4]
  assign mem_0_22_RW0_wmode = RW0_wmode; // @[:anonymous source@296.4]
  assign mem_0_22_RW0_wmask = RW0_wmask[22]; // @[:anonymous source@295.4]
  assign mem_0_23_RW0_addr = RW0_addr; // @[:anonymous source@299.4]
  assign mem_0_23_RW0_clk = RW0_clk; // @[:anonymous source@298.4]
  assign mem_0_23_RW0_wdata = RW0_wdata[191:184]; // @[:anonymous source@301.4]
  assign mem_0_23_RW0_en = RW0_en; // @[:anonymous source@304.4]
  assign mem_0_23_RW0_wmode = RW0_wmode; // @[:anonymous source@303.4]
  assign mem_0_23_RW0_wmask = RW0_wmask[23]; // @[:anonymous source@302.4]
  assign mem_0_24_RW0_addr = RW0_addr; // @[:anonymous source@306.4]
  assign mem_0_24_RW0_clk = RW0_clk; // @[:anonymous source@305.4]
  assign mem_0_24_RW0_wdata = RW0_wdata[199:192]; // @[:anonymous source@308.4]
  assign mem_0_24_RW0_en = RW0_en; // @[:anonymous source@311.4]
  assign mem_0_24_RW0_wmode = RW0_wmode; // @[:anonymous source@310.4]
  assign mem_0_24_RW0_wmask = RW0_wmask[24]; // @[:anonymous source@309.4]
  assign mem_0_25_RW0_addr = RW0_addr; // @[:anonymous source@313.4]
  assign mem_0_25_RW0_clk = RW0_clk; // @[:anonymous source@312.4]
  assign mem_0_25_RW0_wdata = RW0_wdata[207:200]; // @[:anonymous source@315.4]
  assign mem_0_25_RW0_en = RW0_en; // @[:anonymous source@318.4]
  assign mem_0_25_RW0_wmode = RW0_wmode; // @[:anonymous source@317.4]
  assign mem_0_25_RW0_wmask = RW0_wmask[25]; // @[:anonymous source@316.4]
  assign mem_0_26_RW0_addr = RW0_addr; // @[:anonymous source@320.4]
  assign mem_0_26_RW0_clk = RW0_clk; // @[:anonymous source@319.4]
  assign mem_0_26_RW0_wdata = RW0_wdata[215:208]; // @[:anonymous source@322.4]
  assign mem_0_26_RW0_en = RW0_en; // @[:anonymous source@325.4]
  assign mem_0_26_RW0_wmode = RW0_wmode; // @[:anonymous source@324.4]
  assign mem_0_26_RW0_wmask = RW0_wmask[26]; // @[:anonymous source@323.4]
  assign mem_0_27_RW0_addr = RW0_addr; // @[:anonymous source@327.4]
  assign mem_0_27_RW0_clk = RW0_clk; // @[:anonymous source@326.4]
  assign mem_0_27_RW0_wdata = RW0_wdata[223:216]; // @[:anonymous source@329.4]
  assign mem_0_27_RW0_en = RW0_en; // @[:anonymous source@332.4]
  assign mem_0_27_RW0_wmode = RW0_wmode; // @[:anonymous source@331.4]
  assign mem_0_27_RW0_wmask = RW0_wmask[27]; // @[:anonymous source@330.4]
  assign mem_0_28_RW0_addr = RW0_addr; // @[:anonymous source@334.4]
  assign mem_0_28_RW0_clk = RW0_clk; // @[:anonymous source@333.4]
  assign mem_0_28_RW0_wdata = RW0_wdata[231:224]; // @[:anonymous source@336.4]
  assign mem_0_28_RW0_en = RW0_en; // @[:anonymous source@339.4]
  assign mem_0_28_RW0_wmode = RW0_wmode; // @[:anonymous source@338.4]
  assign mem_0_28_RW0_wmask = RW0_wmask[28]; // @[:anonymous source@337.4]
  assign mem_0_29_RW0_addr = RW0_addr; // @[:anonymous source@341.4]
  assign mem_0_29_RW0_clk = RW0_clk; // @[:anonymous source@340.4]
  assign mem_0_29_RW0_wdata = RW0_wdata[239:232]; // @[:anonymous source@343.4]
  assign mem_0_29_RW0_en = RW0_en; // @[:anonymous source@346.4]
  assign mem_0_29_RW0_wmode = RW0_wmode; // @[:anonymous source@345.4]
  assign mem_0_29_RW0_wmask = RW0_wmask[29]; // @[:anonymous source@344.4]
  assign mem_0_30_RW0_addr = RW0_addr; // @[:anonymous source@348.4]
  assign mem_0_30_RW0_clk = RW0_clk; // @[:anonymous source@347.4]
  assign mem_0_30_RW0_wdata = RW0_wdata[247:240]; // @[:anonymous source@350.4]
  assign mem_0_30_RW0_en = RW0_en; // @[:anonymous source@353.4]
  assign mem_0_30_RW0_wmode = RW0_wmode; // @[:anonymous source@352.4]
  assign mem_0_30_RW0_wmask = RW0_wmask[30]; // @[:anonymous source@351.4]
  assign mem_0_31_RW0_addr = RW0_addr; // @[:anonymous source@355.4]
  assign mem_0_31_RW0_clk = RW0_clk; // @[:anonymous source@354.4]
  assign mem_0_31_RW0_wdata = RW0_wdata[255:248]; // @[:anonymous source@357.4]
  assign mem_0_31_RW0_en = RW0_en; // @[:anonymous source@360.4]
  assign mem_0_31_RW0_wmode = RW0_wmode; // @[:anonymous source@359.4]
  assign mem_0_31_RW0_wmask = RW0_wmask[31]; // @[:anonymous source@358.4]
endmodule
module tag_array_ext( // @[:anonymous source@364.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@365.4]
  input         RW0_clk, // @[:anonymous source@366.4]
  input  [87:0] RW0_wdata, // @[:anonymous source@367.4]
  output [87:0] RW0_rdata, // @[:anonymous source@368.4]
  input         RW0_en, // @[:anonymous source@369.4]
  input         RW0_wmode, // @[:anonymous source@370.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@371.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@373.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@373.4]
  wire [21:0] mem_0_0_RW0_wdata; // @[:anonymous source@373.4]
  wire [21:0] mem_0_0_RW0_rdata; // @[:anonymous source@373.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@373.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@373.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@373.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@374.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@374.4]
  wire [21:0] mem_0_1_RW0_wdata; // @[:anonymous source@374.4]
  wire [21:0] mem_0_1_RW0_rdata; // @[:anonymous source@374.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@374.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@374.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@374.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@375.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@375.4]
  wire [21:0] mem_0_2_RW0_wdata; // @[:anonymous source@375.4]
  wire [21:0] mem_0_2_RW0_rdata; // @[:anonymous source@375.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@375.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@375.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@375.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@376.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@376.4]
  wire [21:0] mem_0_3_RW0_wdata; // @[:anonymous source@376.4]
  wire [21:0] mem_0_3_RW0_rdata; // @[:anonymous source@376.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@376.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@376.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@376.4]
  wire [21:0] RW0_rdata_0_0; // @[:anonymous source@379.4]
  wire [21:0] RW0_rdata_0_1; // @[:anonymous source@386.4]
  wire [21:0] RW0_rdata_0_2; // @[:anonymous source@393.4]
  wire [21:0] RW0_rdata_0_3; // @[:anonymous source@400.4]
  wire [43:0] _GEN_0; // @[:anonymous source@405.4]
  wire [65:0] _GEN_1; // @[:anonymous source@405.4]
  wire [87:0] RW0_rdata_0; // @[:anonymous source@405.4]
  wire [43:0] _GEN_2; // @[:anonymous source@406.4]
  wire [65:0] _GEN_3; // @[:anonymous source@406.4]
  split_tag_array_ext mem_0_0 ( // @[:anonymous source@373.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 ( // @[:anonymous source@374.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 ( // @[:anonymous source@375.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 ( // @[:anonymous source@376.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@379.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@386.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@393.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@400.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@405.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@405.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@405.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@406.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@406.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@406.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@378.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@377.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0]; // @[:anonymous source@380.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@383.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@382.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@381.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@385.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@384.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22]; // @[:anonymous source@387.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@390.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@389.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@388.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@392.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@391.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44]; // @[:anonymous source@394.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@397.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@396.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@395.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@399.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@398.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66]; // @[:anonymous source@401.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@404.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@403.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@402.4]
endmodule
module mem_ext( // @[:anonymous source@408.2]
  input  [11:0]  W0_addr, // @[:anonymous source@409.4]
  input          W0_clk, // @[:anonymous source@410.4]
  input  [127:0] W0_data, // @[:anonymous source@411.4]
  input          W0_en, // @[:anonymous source@412.4]
  input  [15:0]  W0_mask, // @[:anonymous source@413.4]
  input  [11:0]  R0_addr, // @[:anonymous source@414.4]
  input          R0_clk, // @[:anonymous source@415.4]
  output [127:0] R0_data, // @[:anonymous source@416.4]
  input          R0_en // @[:anonymous source@417.4]
);
  wire [11:0] mem_0_0_W0_addr; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@419.4]
  wire [7:0] mem_0_0_W0_data; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@419.4]
  wire [11:0] mem_0_0_R0_addr; // @[:anonymous source@419.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@419.4]
  wire [7:0] mem_0_0_R0_data; // @[:anonymous source@419.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@419.4]
  wire [11:0] mem_0_1_W0_addr; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@420.4]
  wire [7:0] mem_0_1_W0_data; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@420.4]
  wire [11:0] mem_0_1_R0_addr; // @[:anonymous source@420.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@420.4]
  wire [7:0] mem_0_1_R0_data; // @[:anonymous source@420.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@420.4]
  wire [11:0] mem_0_2_W0_addr; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@421.4]
  wire [7:0] mem_0_2_W0_data; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@421.4]
  wire [11:0] mem_0_2_R0_addr; // @[:anonymous source@421.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@421.4]
  wire [7:0] mem_0_2_R0_data; // @[:anonymous source@421.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@421.4]
  wire [11:0] mem_0_3_W0_addr; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@422.4]
  wire [7:0] mem_0_3_W0_data; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@422.4]
  wire [11:0] mem_0_3_R0_addr; // @[:anonymous source@422.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@422.4]
  wire [7:0] mem_0_3_R0_data; // @[:anonymous source@422.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@422.4]
  wire [11:0] mem_0_4_W0_addr; // @[:anonymous source@423.4]
  wire  mem_0_4_W0_clk; // @[:anonymous source@423.4]
  wire [7:0] mem_0_4_W0_data; // @[:anonymous source@423.4]
  wire  mem_0_4_W0_en; // @[:anonymous source@423.4]
  wire  mem_0_4_W0_mask; // @[:anonymous source@423.4]
  wire [11:0] mem_0_4_R0_addr; // @[:anonymous source@423.4]
  wire  mem_0_4_R0_clk; // @[:anonymous source@423.4]
  wire [7:0] mem_0_4_R0_data; // @[:anonymous source@423.4]
  wire  mem_0_4_R0_en; // @[:anonymous source@423.4]
  wire [11:0] mem_0_5_W0_addr; // @[:anonymous source@424.4]
  wire  mem_0_5_W0_clk; // @[:anonymous source@424.4]
  wire [7:0] mem_0_5_W0_data; // @[:anonymous source@424.4]
  wire  mem_0_5_W0_en; // @[:anonymous source@424.4]
  wire  mem_0_5_W0_mask; // @[:anonymous source@424.4]
  wire [11:0] mem_0_5_R0_addr; // @[:anonymous source@424.4]
  wire  mem_0_5_R0_clk; // @[:anonymous source@424.4]
  wire [7:0] mem_0_5_R0_data; // @[:anonymous source@424.4]
  wire  mem_0_5_R0_en; // @[:anonymous source@424.4]
  wire [11:0] mem_0_6_W0_addr; // @[:anonymous source@425.4]
  wire  mem_0_6_W0_clk; // @[:anonymous source@425.4]
  wire [7:0] mem_0_6_W0_data; // @[:anonymous source@425.4]
  wire  mem_0_6_W0_en; // @[:anonymous source@425.4]
  wire  mem_0_6_W0_mask; // @[:anonymous source@425.4]
  wire [11:0] mem_0_6_R0_addr; // @[:anonymous source@425.4]
  wire  mem_0_6_R0_clk; // @[:anonymous source@425.4]
  wire [7:0] mem_0_6_R0_data; // @[:anonymous source@425.4]
  wire  mem_0_6_R0_en; // @[:anonymous source@425.4]
  wire [11:0] mem_0_7_W0_addr; // @[:anonymous source@426.4]
  wire  mem_0_7_W0_clk; // @[:anonymous source@426.4]
  wire [7:0] mem_0_7_W0_data; // @[:anonymous source@426.4]
  wire  mem_0_7_W0_en; // @[:anonymous source@426.4]
  wire  mem_0_7_W0_mask; // @[:anonymous source@426.4]
  wire [11:0] mem_0_7_R0_addr; // @[:anonymous source@426.4]
  wire  mem_0_7_R0_clk; // @[:anonymous source@426.4]
  wire [7:0] mem_0_7_R0_data; // @[:anonymous source@426.4]
  wire  mem_0_7_R0_en; // @[:anonymous source@426.4]
  wire [11:0] mem_0_8_W0_addr; // @[:anonymous source@427.4]
  wire  mem_0_8_W0_clk; // @[:anonymous source@427.4]
  wire [7:0] mem_0_8_W0_data; // @[:anonymous source@427.4]
  wire  mem_0_8_W0_en; // @[:anonymous source@427.4]
  wire  mem_0_8_W0_mask; // @[:anonymous source@427.4]
  wire [11:0] mem_0_8_R0_addr; // @[:anonymous source@427.4]
  wire  mem_0_8_R0_clk; // @[:anonymous source@427.4]
  wire [7:0] mem_0_8_R0_data; // @[:anonymous source@427.4]
  wire  mem_0_8_R0_en; // @[:anonymous source@427.4]
  wire [11:0] mem_0_9_W0_addr; // @[:anonymous source@428.4]
  wire  mem_0_9_W0_clk; // @[:anonymous source@428.4]
  wire [7:0] mem_0_9_W0_data; // @[:anonymous source@428.4]
  wire  mem_0_9_W0_en; // @[:anonymous source@428.4]
  wire  mem_0_9_W0_mask; // @[:anonymous source@428.4]
  wire [11:0] mem_0_9_R0_addr; // @[:anonymous source@428.4]
  wire  mem_0_9_R0_clk; // @[:anonymous source@428.4]
  wire [7:0] mem_0_9_R0_data; // @[:anonymous source@428.4]
  wire  mem_0_9_R0_en; // @[:anonymous source@428.4]
  wire [11:0] mem_0_10_W0_addr; // @[:anonymous source@429.4]
  wire  mem_0_10_W0_clk; // @[:anonymous source@429.4]
  wire [7:0] mem_0_10_W0_data; // @[:anonymous source@429.4]
  wire  mem_0_10_W0_en; // @[:anonymous source@429.4]
  wire  mem_0_10_W0_mask; // @[:anonymous source@429.4]
  wire [11:0] mem_0_10_R0_addr; // @[:anonymous source@429.4]
  wire  mem_0_10_R0_clk; // @[:anonymous source@429.4]
  wire [7:0] mem_0_10_R0_data; // @[:anonymous source@429.4]
  wire  mem_0_10_R0_en; // @[:anonymous source@429.4]
  wire [11:0] mem_0_11_W0_addr; // @[:anonymous source@430.4]
  wire  mem_0_11_W0_clk; // @[:anonymous source@430.4]
  wire [7:0] mem_0_11_W0_data; // @[:anonymous source@430.4]
  wire  mem_0_11_W0_en; // @[:anonymous source@430.4]
  wire  mem_0_11_W0_mask; // @[:anonymous source@430.4]
  wire [11:0] mem_0_11_R0_addr; // @[:anonymous source@430.4]
  wire  mem_0_11_R0_clk; // @[:anonymous source@430.4]
  wire [7:0] mem_0_11_R0_data; // @[:anonymous source@430.4]
  wire  mem_0_11_R0_en; // @[:anonymous source@430.4]
  wire [11:0] mem_0_12_W0_addr; // @[:anonymous source@431.4]
  wire  mem_0_12_W0_clk; // @[:anonymous source@431.4]
  wire [7:0] mem_0_12_W0_data; // @[:anonymous source@431.4]
  wire  mem_0_12_W0_en; // @[:anonymous source@431.4]
  wire  mem_0_12_W0_mask; // @[:anonymous source@431.4]
  wire [11:0] mem_0_12_R0_addr; // @[:anonymous source@431.4]
  wire  mem_0_12_R0_clk; // @[:anonymous source@431.4]
  wire [7:0] mem_0_12_R0_data; // @[:anonymous source@431.4]
  wire  mem_0_12_R0_en; // @[:anonymous source@431.4]
  wire [11:0] mem_0_13_W0_addr; // @[:anonymous source@432.4]
  wire  mem_0_13_W0_clk; // @[:anonymous source@432.4]
  wire [7:0] mem_0_13_W0_data; // @[:anonymous source@432.4]
  wire  mem_0_13_W0_en; // @[:anonymous source@432.4]
  wire  mem_0_13_W0_mask; // @[:anonymous source@432.4]
  wire [11:0] mem_0_13_R0_addr; // @[:anonymous source@432.4]
  wire  mem_0_13_R0_clk; // @[:anonymous source@432.4]
  wire [7:0] mem_0_13_R0_data; // @[:anonymous source@432.4]
  wire  mem_0_13_R0_en; // @[:anonymous source@432.4]
  wire [11:0] mem_0_14_W0_addr; // @[:anonymous source@433.4]
  wire  mem_0_14_W0_clk; // @[:anonymous source@433.4]
  wire [7:0] mem_0_14_W0_data; // @[:anonymous source@433.4]
  wire  mem_0_14_W0_en; // @[:anonymous source@433.4]
  wire  mem_0_14_W0_mask; // @[:anonymous source@433.4]
  wire [11:0] mem_0_14_R0_addr; // @[:anonymous source@433.4]
  wire  mem_0_14_R0_clk; // @[:anonymous source@433.4]
  wire [7:0] mem_0_14_R0_data; // @[:anonymous source@433.4]
  wire  mem_0_14_R0_en; // @[:anonymous source@433.4]
  wire [11:0] mem_0_15_W0_addr; // @[:anonymous source@434.4]
  wire  mem_0_15_W0_clk; // @[:anonymous source@434.4]
  wire [7:0] mem_0_15_W0_data; // @[:anonymous source@434.4]
  wire  mem_0_15_W0_en; // @[:anonymous source@434.4]
  wire  mem_0_15_W0_mask; // @[:anonymous source@434.4]
  wire [11:0] mem_0_15_R0_addr; // @[:anonymous source@434.4]
  wire  mem_0_15_R0_clk; // @[:anonymous source@434.4]
  wire [7:0] mem_0_15_R0_data; // @[:anonymous source@434.4]
  wire  mem_0_15_R0_en; // @[:anonymous source@434.4]
  wire [7:0] R0_data_0_0; // @[:anonymous source@517.4]
  wire [7:0] R0_data_0_1; // @[:anonymous source@521.4]
  wire [7:0] R0_data_0_2; // @[:anonymous source@525.4]
  wire [7:0] R0_data_0_3; // @[:anonymous source@529.4]
  wire [7:0] R0_data_0_4; // @[:anonymous source@533.4]
  wire [7:0] R0_data_0_5; // @[:anonymous source@537.4]
  wire [7:0] R0_data_0_6; // @[:anonymous source@541.4]
  wire [7:0] R0_data_0_7; // @[:anonymous source@545.4]
  wire [7:0] R0_data_0_8; // @[:anonymous source@549.4]
  wire [7:0] R0_data_0_9; // @[:anonymous source@553.4]
  wire [7:0] R0_data_0_10; // @[:anonymous source@557.4]
  wire [7:0] R0_data_0_11; // @[:anonymous source@561.4]
  wire [7:0] R0_data_0_12; // @[:anonymous source@565.4]
  wire [7:0] R0_data_0_13; // @[:anonymous source@569.4]
  wire [7:0] R0_data_0_14; // @[:anonymous source@573.4]
  wire [7:0] R0_data_0_15; // @[:anonymous source@577.4]
  wire [15:0] _GEN_0; // @[:anonymous source@579.4]
  wire [23:0] _GEN_1; // @[:anonymous source@579.4]
  wire [31:0] _GEN_2; // @[:anonymous source@579.4]
  wire [39:0] _GEN_3; // @[:anonymous source@579.4]
  wire [47:0] _GEN_4; // @[:anonymous source@579.4]
  wire [55:0] _GEN_5; // @[:anonymous source@579.4]
  wire [63:0] _GEN_6; // @[:anonymous source@579.4]
  wire [71:0] _GEN_7; // @[:anonymous source@579.4]
  wire [79:0] _GEN_8; // @[:anonymous source@579.4]
  wire [87:0] _GEN_9; // @[:anonymous source@579.4]
  wire [95:0] _GEN_10; // @[:anonymous source@579.4]
  wire [103:0] _GEN_11; // @[:anonymous source@579.4]
  wire [111:0] _GEN_12; // @[:anonymous source@579.4]
  wire [119:0] _GEN_13; // @[:anonymous source@579.4]
  wire [127:0] R0_data_0; // @[:anonymous source@579.4]
  wire [15:0] _GEN_14; // @[:anonymous source@580.4]
  wire [23:0] _GEN_15; // @[:anonymous source@580.4]
  wire [31:0] _GEN_16; // @[:anonymous source@580.4]
  wire [39:0] _GEN_17; // @[:anonymous source@580.4]
  wire [47:0] _GEN_18; // @[:anonymous source@580.4]
  wire [55:0] _GEN_19; // @[:anonymous source@580.4]
  wire [63:0] _GEN_20; // @[:anonymous source@580.4]
  wire [71:0] _GEN_21; // @[:anonymous source@580.4]
  wire [79:0] _GEN_22; // @[:anonymous source@580.4]
  wire [87:0] _GEN_23; // @[:anonymous source@580.4]
  wire [95:0] _GEN_24; // @[:anonymous source@580.4]
  wire [103:0] _GEN_25; // @[:anonymous source@580.4]
  wire [111:0] _GEN_26; // @[:anonymous source@580.4]
  wire [119:0] _GEN_27; // @[:anonymous source@580.4]
  split_mem_ext mem_0_0 ( // @[:anonymous source@419.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_mem_ext mem_0_1 ( // @[:anonymous source@420.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_mem_ext mem_0_2 ( // @[:anonymous source@421.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_mem_ext mem_0_3 ( // @[:anonymous source@422.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  split_mem_ext mem_0_4 ( // @[:anonymous source@423.4]
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask),
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en)
  );
  split_mem_ext mem_0_5 ( // @[:anonymous source@424.4]
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask),
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en)
  );
  split_mem_ext mem_0_6 ( // @[:anonymous source@425.4]
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask),
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en)
  );
  split_mem_ext mem_0_7 ( // @[:anonymous source@426.4]
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask),
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en)
  );
  split_mem_ext mem_0_8 ( // @[:anonymous source@427.4]
    .W0_addr(mem_0_8_W0_addr),
    .W0_clk(mem_0_8_W0_clk),
    .W0_data(mem_0_8_W0_data),
    .W0_en(mem_0_8_W0_en),
    .W0_mask(mem_0_8_W0_mask),
    .R0_addr(mem_0_8_R0_addr),
    .R0_clk(mem_0_8_R0_clk),
    .R0_data(mem_0_8_R0_data),
    .R0_en(mem_0_8_R0_en)
  );
  split_mem_ext mem_0_9 ( // @[:anonymous source@428.4]
    .W0_addr(mem_0_9_W0_addr),
    .W0_clk(mem_0_9_W0_clk),
    .W0_data(mem_0_9_W0_data),
    .W0_en(mem_0_9_W0_en),
    .W0_mask(mem_0_9_W0_mask),
    .R0_addr(mem_0_9_R0_addr),
    .R0_clk(mem_0_9_R0_clk),
    .R0_data(mem_0_9_R0_data),
    .R0_en(mem_0_9_R0_en)
  );
  split_mem_ext mem_0_10 ( // @[:anonymous source@429.4]
    .W0_addr(mem_0_10_W0_addr),
    .W0_clk(mem_0_10_W0_clk),
    .W0_data(mem_0_10_W0_data),
    .W0_en(mem_0_10_W0_en),
    .W0_mask(mem_0_10_W0_mask),
    .R0_addr(mem_0_10_R0_addr),
    .R0_clk(mem_0_10_R0_clk),
    .R0_data(mem_0_10_R0_data),
    .R0_en(mem_0_10_R0_en)
  );
  split_mem_ext mem_0_11 ( // @[:anonymous source@430.4]
    .W0_addr(mem_0_11_W0_addr),
    .W0_clk(mem_0_11_W0_clk),
    .W0_data(mem_0_11_W0_data),
    .W0_en(mem_0_11_W0_en),
    .W0_mask(mem_0_11_W0_mask),
    .R0_addr(mem_0_11_R0_addr),
    .R0_clk(mem_0_11_R0_clk),
    .R0_data(mem_0_11_R0_data),
    .R0_en(mem_0_11_R0_en)
  );
  split_mem_ext mem_0_12 ( // @[:anonymous source@431.4]
    .W0_addr(mem_0_12_W0_addr),
    .W0_clk(mem_0_12_W0_clk),
    .W0_data(mem_0_12_W0_data),
    .W0_en(mem_0_12_W0_en),
    .W0_mask(mem_0_12_W0_mask),
    .R0_addr(mem_0_12_R0_addr),
    .R0_clk(mem_0_12_R0_clk),
    .R0_data(mem_0_12_R0_data),
    .R0_en(mem_0_12_R0_en)
  );
  split_mem_ext mem_0_13 ( // @[:anonymous source@432.4]
    .W0_addr(mem_0_13_W0_addr),
    .W0_clk(mem_0_13_W0_clk),
    .W0_data(mem_0_13_W0_data),
    .W0_en(mem_0_13_W0_en),
    .W0_mask(mem_0_13_W0_mask),
    .R0_addr(mem_0_13_R0_addr),
    .R0_clk(mem_0_13_R0_clk),
    .R0_data(mem_0_13_R0_data),
    .R0_en(mem_0_13_R0_en)
  );
  split_mem_ext mem_0_14 ( // @[:anonymous source@433.4]
    .W0_addr(mem_0_14_W0_addr),
    .W0_clk(mem_0_14_W0_clk),
    .W0_data(mem_0_14_W0_data),
    .W0_en(mem_0_14_W0_en),
    .W0_mask(mem_0_14_W0_mask),
    .R0_addr(mem_0_14_R0_addr),
    .R0_clk(mem_0_14_R0_clk),
    .R0_data(mem_0_14_R0_data),
    .R0_en(mem_0_14_R0_en)
  );
  split_mem_ext mem_0_15 ( // @[:anonymous source@434.4]
    .W0_addr(mem_0_15_W0_addr),
    .W0_clk(mem_0_15_W0_clk),
    .W0_data(mem_0_15_W0_data),
    .W0_en(mem_0_15_W0_en),
    .W0_mask(mem_0_15_W0_mask),
    .R0_addr(mem_0_15_R0_addr),
    .R0_clk(mem_0_15_R0_clk),
    .R0_data(mem_0_15_R0_data),
    .R0_en(mem_0_15_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@517.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@521.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@525.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@529.4]
  assign R0_data_0_4 = mem_0_4_R0_data; // @[:anonymous source@533.4]
  assign R0_data_0_5 = mem_0_5_R0_data; // @[:anonymous source@537.4]
  assign R0_data_0_6 = mem_0_6_R0_data; // @[:anonymous source@541.4]
  assign R0_data_0_7 = mem_0_7_R0_data; // @[:anonymous source@545.4]
  assign R0_data_0_8 = mem_0_8_R0_data; // @[:anonymous source@549.4]
  assign R0_data_0_9 = mem_0_9_R0_data; // @[:anonymous source@553.4]
  assign R0_data_0_10 = mem_0_10_R0_data; // @[:anonymous source@557.4]
  assign R0_data_0_11 = mem_0_11_R0_data; // @[:anonymous source@561.4]
  assign R0_data_0_12 = mem_0_12_R0_data; // @[:anonymous source@565.4]
  assign R0_data_0_13 = mem_0_13_R0_data; // @[:anonymous source@569.4]
  assign R0_data_0_14 = mem_0_14_R0_data; // @[:anonymous source@573.4]
  assign R0_data_0_15 = mem_0_15_R0_data; // @[:anonymous source@577.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_2 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_3 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_4 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_5 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_6 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_7 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_8 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@579.4]
  assign _GEN_9 = {R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign _GEN_10 = {R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign _GEN_11 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign _GEN_12 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign _GEN_13 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign R0_data_0 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@579.4]
  assign _GEN_14 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_15 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_16 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_17 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_18 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_19 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_20 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_21 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_22 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@580.4]
  assign _GEN_23 = {R0_data_0_10,_GEN_8}; // @[:anonymous source@580.4]
  assign _GEN_24 = {R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@580.4]
  assign _GEN_25 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@580.4]
  assign _GEN_26 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@580.4]
  assign _GEN_27 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@580.4]
  assign R0_data = {R0_data_0_15,_GEN_13}; // @[:anonymous source@580.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@436.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@435.4]
  assign mem_0_0_W0_data = W0_data[7:0]; // @[:anonymous source@437.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@439.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@438.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@516.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@515.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@518.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@441.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@440.4]
  assign mem_0_1_W0_data = W0_data[15:8]; // @[:anonymous source@442.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@444.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@443.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@520.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@519.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@522.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@446.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@445.4]
  assign mem_0_2_W0_data = W0_data[23:16]; // @[:anonymous source@447.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@449.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@448.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@524.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@523.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@526.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@451.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@450.4]
  assign mem_0_3_W0_data = W0_data[31:24]; // @[:anonymous source@452.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@454.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@453.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@528.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@527.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@530.4]
  assign mem_0_4_W0_addr = W0_addr; // @[:anonymous source@456.4]
  assign mem_0_4_W0_clk = W0_clk; // @[:anonymous source@455.4]
  assign mem_0_4_W0_data = W0_data[39:32]; // @[:anonymous source@457.4]
  assign mem_0_4_W0_en = W0_en; // @[:anonymous source@459.4]
  assign mem_0_4_W0_mask = W0_mask[4]; // @[:anonymous source@458.4]
  assign mem_0_4_R0_addr = R0_addr; // @[:anonymous source@532.4]
  assign mem_0_4_R0_clk = R0_clk; // @[:anonymous source@531.4]
  assign mem_0_4_R0_en = R0_en; // @[:anonymous source@534.4]
  assign mem_0_5_W0_addr = W0_addr; // @[:anonymous source@461.4]
  assign mem_0_5_W0_clk = W0_clk; // @[:anonymous source@460.4]
  assign mem_0_5_W0_data = W0_data[47:40]; // @[:anonymous source@462.4]
  assign mem_0_5_W0_en = W0_en; // @[:anonymous source@464.4]
  assign mem_0_5_W0_mask = W0_mask[5]; // @[:anonymous source@463.4]
  assign mem_0_5_R0_addr = R0_addr; // @[:anonymous source@536.4]
  assign mem_0_5_R0_clk = R0_clk; // @[:anonymous source@535.4]
  assign mem_0_5_R0_en = R0_en; // @[:anonymous source@538.4]
  assign mem_0_6_W0_addr = W0_addr; // @[:anonymous source@466.4]
  assign mem_0_6_W0_clk = W0_clk; // @[:anonymous source@465.4]
  assign mem_0_6_W0_data = W0_data[55:48]; // @[:anonymous source@467.4]
  assign mem_0_6_W0_en = W0_en; // @[:anonymous source@469.4]
  assign mem_0_6_W0_mask = W0_mask[6]; // @[:anonymous source@468.4]
  assign mem_0_6_R0_addr = R0_addr; // @[:anonymous source@540.4]
  assign mem_0_6_R0_clk = R0_clk; // @[:anonymous source@539.4]
  assign mem_0_6_R0_en = R0_en; // @[:anonymous source@542.4]
  assign mem_0_7_W0_addr = W0_addr; // @[:anonymous source@471.4]
  assign mem_0_7_W0_clk = W0_clk; // @[:anonymous source@470.4]
  assign mem_0_7_W0_data = W0_data[63:56]; // @[:anonymous source@472.4]
  assign mem_0_7_W0_en = W0_en; // @[:anonymous source@474.4]
  assign mem_0_7_W0_mask = W0_mask[7]; // @[:anonymous source@473.4]
  assign mem_0_7_R0_addr = R0_addr; // @[:anonymous source@544.4]
  assign mem_0_7_R0_clk = R0_clk; // @[:anonymous source@543.4]
  assign mem_0_7_R0_en = R0_en; // @[:anonymous source@546.4]
  assign mem_0_8_W0_addr = W0_addr; // @[:anonymous source@476.4]
  assign mem_0_8_W0_clk = W0_clk; // @[:anonymous source@475.4]
  assign mem_0_8_W0_data = W0_data[71:64]; // @[:anonymous source@477.4]
  assign mem_0_8_W0_en = W0_en; // @[:anonymous source@479.4]
  assign mem_0_8_W0_mask = W0_mask[8]; // @[:anonymous source@478.4]
  assign mem_0_8_R0_addr = R0_addr; // @[:anonymous source@548.4]
  assign mem_0_8_R0_clk = R0_clk; // @[:anonymous source@547.4]
  assign mem_0_8_R0_en = R0_en; // @[:anonymous source@550.4]
  assign mem_0_9_W0_addr = W0_addr; // @[:anonymous source@481.4]
  assign mem_0_9_W0_clk = W0_clk; // @[:anonymous source@480.4]
  assign mem_0_9_W0_data = W0_data[79:72]; // @[:anonymous source@482.4]
  assign mem_0_9_W0_en = W0_en; // @[:anonymous source@484.4]
  assign mem_0_9_W0_mask = W0_mask[9]; // @[:anonymous source@483.4]
  assign mem_0_9_R0_addr = R0_addr; // @[:anonymous source@552.4]
  assign mem_0_9_R0_clk = R0_clk; // @[:anonymous source@551.4]
  assign mem_0_9_R0_en = R0_en; // @[:anonymous source@554.4]
  assign mem_0_10_W0_addr = W0_addr; // @[:anonymous source@486.4]
  assign mem_0_10_W0_clk = W0_clk; // @[:anonymous source@485.4]
  assign mem_0_10_W0_data = W0_data[87:80]; // @[:anonymous source@487.4]
  assign mem_0_10_W0_en = W0_en; // @[:anonymous source@489.4]
  assign mem_0_10_W0_mask = W0_mask[10]; // @[:anonymous source@488.4]
  assign mem_0_10_R0_addr = R0_addr; // @[:anonymous source@556.4]
  assign mem_0_10_R0_clk = R0_clk; // @[:anonymous source@555.4]
  assign mem_0_10_R0_en = R0_en; // @[:anonymous source@558.4]
  assign mem_0_11_W0_addr = W0_addr; // @[:anonymous source@491.4]
  assign mem_0_11_W0_clk = W0_clk; // @[:anonymous source@490.4]
  assign mem_0_11_W0_data = W0_data[95:88]; // @[:anonymous source@492.4]
  assign mem_0_11_W0_en = W0_en; // @[:anonymous source@494.4]
  assign mem_0_11_W0_mask = W0_mask[11]; // @[:anonymous source@493.4]
  assign mem_0_11_R0_addr = R0_addr; // @[:anonymous source@560.4]
  assign mem_0_11_R0_clk = R0_clk; // @[:anonymous source@559.4]
  assign mem_0_11_R0_en = R0_en; // @[:anonymous source@562.4]
  assign mem_0_12_W0_addr = W0_addr; // @[:anonymous source@496.4]
  assign mem_0_12_W0_clk = W0_clk; // @[:anonymous source@495.4]
  assign mem_0_12_W0_data = W0_data[103:96]; // @[:anonymous source@497.4]
  assign mem_0_12_W0_en = W0_en; // @[:anonymous source@499.4]
  assign mem_0_12_W0_mask = W0_mask[12]; // @[:anonymous source@498.4]
  assign mem_0_12_R0_addr = R0_addr; // @[:anonymous source@564.4]
  assign mem_0_12_R0_clk = R0_clk; // @[:anonymous source@563.4]
  assign mem_0_12_R0_en = R0_en; // @[:anonymous source@566.4]
  assign mem_0_13_W0_addr = W0_addr; // @[:anonymous source@501.4]
  assign mem_0_13_W0_clk = W0_clk; // @[:anonymous source@500.4]
  assign mem_0_13_W0_data = W0_data[111:104]; // @[:anonymous source@502.4]
  assign mem_0_13_W0_en = W0_en; // @[:anonymous source@504.4]
  assign mem_0_13_W0_mask = W0_mask[13]; // @[:anonymous source@503.4]
  assign mem_0_13_R0_addr = R0_addr; // @[:anonymous source@568.4]
  assign mem_0_13_R0_clk = R0_clk; // @[:anonymous source@567.4]
  assign mem_0_13_R0_en = R0_en; // @[:anonymous source@570.4]
  assign mem_0_14_W0_addr = W0_addr; // @[:anonymous source@506.4]
  assign mem_0_14_W0_clk = W0_clk; // @[:anonymous source@505.4]
  assign mem_0_14_W0_data = W0_data[119:112]; // @[:anonymous source@507.4]
  assign mem_0_14_W0_en = W0_en; // @[:anonymous source@509.4]
  assign mem_0_14_W0_mask = W0_mask[14]; // @[:anonymous source@508.4]
  assign mem_0_14_R0_addr = R0_addr; // @[:anonymous source@572.4]
  assign mem_0_14_R0_clk = R0_clk; // @[:anonymous source@571.4]
  assign mem_0_14_R0_en = R0_en; // @[:anonymous source@574.4]
  assign mem_0_15_W0_addr = W0_addr; // @[:anonymous source@511.4]
  assign mem_0_15_W0_clk = W0_clk; // @[:anonymous source@510.4]
  assign mem_0_15_W0_data = W0_data[127:120]; // @[:anonymous source@512.4]
  assign mem_0_15_W0_en = W0_en; // @[:anonymous source@514.4]
  assign mem_0_15_W0_mask = W0_mask[15]; // @[:anonymous source@513.4]
  assign mem_0_15_R0_addr = R0_addr; // @[:anonymous source@576.4]
  assign mem_0_15_R0_clk = R0_clk; // @[:anonymous source@575.4]
  assign mem_0_15_R0_en = R0_en; // @[:anonymous source@578.4]
endmodule
module mem_0_ext( // @[:anonymous source@582.2]
  input  [9:0]   W0_addr, // @[:anonymous source@583.4]
  input          W0_clk, // @[:anonymous source@584.4]
  input  [511:0] W0_data, // @[:anonymous source@585.4]
  input          W0_en, // @[:anonymous source@586.4]
  input  [63:0]  W0_mask, // @[:anonymous source@587.4]
  input  [9:0]   R0_addr, // @[:anonymous source@588.4]
  input          R0_clk, // @[:anonymous source@589.4]
  output [511:0] R0_data, // @[:anonymous source@590.4]
  input          R0_en // @[:anonymous source@591.4]
);
  wire [9:0] mem_0_0_W0_addr; // @[:anonymous source@593.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@593.4]
  wire [7:0] mem_0_0_W0_data; // @[:anonymous source@593.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@593.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@593.4]
  wire [9:0] mem_0_0_R0_addr; // @[:anonymous source@593.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@593.4]
  wire [7:0] mem_0_0_R0_data; // @[:anonymous source@593.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@593.4]
  wire [9:0] mem_0_1_W0_addr; // @[:anonymous source@594.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@594.4]
  wire [7:0] mem_0_1_W0_data; // @[:anonymous source@594.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@594.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@594.4]
  wire [9:0] mem_0_1_R0_addr; // @[:anonymous source@594.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@594.4]
  wire [7:0] mem_0_1_R0_data; // @[:anonymous source@594.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@594.4]
  wire [9:0] mem_0_2_W0_addr; // @[:anonymous source@595.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@595.4]
  wire [7:0] mem_0_2_W0_data; // @[:anonymous source@595.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@595.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@595.4]
  wire [9:0] mem_0_2_R0_addr; // @[:anonymous source@595.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@595.4]
  wire [7:0] mem_0_2_R0_data; // @[:anonymous source@595.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@595.4]
  wire [9:0] mem_0_3_W0_addr; // @[:anonymous source@596.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@596.4]
  wire [7:0] mem_0_3_W0_data; // @[:anonymous source@596.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@596.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@596.4]
  wire [9:0] mem_0_3_R0_addr; // @[:anonymous source@596.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@596.4]
  wire [7:0] mem_0_3_R0_data; // @[:anonymous source@596.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@596.4]
  wire [9:0] mem_0_4_W0_addr; // @[:anonymous source@597.4]
  wire  mem_0_4_W0_clk; // @[:anonymous source@597.4]
  wire [7:0] mem_0_4_W0_data; // @[:anonymous source@597.4]
  wire  mem_0_4_W0_en; // @[:anonymous source@597.4]
  wire  mem_0_4_W0_mask; // @[:anonymous source@597.4]
  wire [9:0] mem_0_4_R0_addr; // @[:anonymous source@597.4]
  wire  mem_0_4_R0_clk; // @[:anonymous source@597.4]
  wire [7:0] mem_0_4_R0_data; // @[:anonymous source@597.4]
  wire  mem_0_4_R0_en; // @[:anonymous source@597.4]
  wire [9:0] mem_0_5_W0_addr; // @[:anonymous source@598.4]
  wire  mem_0_5_W0_clk; // @[:anonymous source@598.4]
  wire [7:0] mem_0_5_W0_data; // @[:anonymous source@598.4]
  wire  mem_0_5_W0_en; // @[:anonymous source@598.4]
  wire  mem_0_5_W0_mask; // @[:anonymous source@598.4]
  wire [9:0] mem_0_5_R0_addr; // @[:anonymous source@598.4]
  wire  mem_0_5_R0_clk; // @[:anonymous source@598.4]
  wire [7:0] mem_0_5_R0_data; // @[:anonymous source@598.4]
  wire  mem_0_5_R0_en; // @[:anonymous source@598.4]
  wire [9:0] mem_0_6_W0_addr; // @[:anonymous source@599.4]
  wire  mem_0_6_W0_clk; // @[:anonymous source@599.4]
  wire [7:0] mem_0_6_W0_data; // @[:anonymous source@599.4]
  wire  mem_0_6_W0_en; // @[:anonymous source@599.4]
  wire  mem_0_6_W0_mask; // @[:anonymous source@599.4]
  wire [9:0] mem_0_6_R0_addr; // @[:anonymous source@599.4]
  wire  mem_0_6_R0_clk; // @[:anonymous source@599.4]
  wire [7:0] mem_0_6_R0_data; // @[:anonymous source@599.4]
  wire  mem_0_6_R0_en; // @[:anonymous source@599.4]
  wire [9:0] mem_0_7_W0_addr; // @[:anonymous source@600.4]
  wire  mem_0_7_W0_clk; // @[:anonymous source@600.4]
  wire [7:0] mem_0_7_W0_data; // @[:anonymous source@600.4]
  wire  mem_0_7_W0_en; // @[:anonymous source@600.4]
  wire  mem_0_7_W0_mask; // @[:anonymous source@600.4]
  wire [9:0] mem_0_7_R0_addr; // @[:anonymous source@600.4]
  wire  mem_0_7_R0_clk; // @[:anonymous source@600.4]
  wire [7:0] mem_0_7_R0_data; // @[:anonymous source@600.4]
  wire  mem_0_7_R0_en; // @[:anonymous source@600.4]
  wire [9:0] mem_0_8_W0_addr; // @[:anonymous source@601.4]
  wire  mem_0_8_W0_clk; // @[:anonymous source@601.4]
  wire [7:0] mem_0_8_W0_data; // @[:anonymous source@601.4]
  wire  mem_0_8_W0_en; // @[:anonymous source@601.4]
  wire  mem_0_8_W0_mask; // @[:anonymous source@601.4]
  wire [9:0] mem_0_8_R0_addr; // @[:anonymous source@601.4]
  wire  mem_0_8_R0_clk; // @[:anonymous source@601.4]
  wire [7:0] mem_0_8_R0_data; // @[:anonymous source@601.4]
  wire  mem_0_8_R0_en; // @[:anonymous source@601.4]
  wire [9:0] mem_0_9_W0_addr; // @[:anonymous source@602.4]
  wire  mem_0_9_W0_clk; // @[:anonymous source@602.4]
  wire [7:0] mem_0_9_W0_data; // @[:anonymous source@602.4]
  wire  mem_0_9_W0_en; // @[:anonymous source@602.4]
  wire  mem_0_9_W0_mask; // @[:anonymous source@602.4]
  wire [9:0] mem_0_9_R0_addr; // @[:anonymous source@602.4]
  wire  mem_0_9_R0_clk; // @[:anonymous source@602.4]
  wire [7:0] mem_0_9_R0_data; // @[:anonymous source@602.4]
  wire  mem_0_9_R0_en; // @[:anonymous source@602.4]
  wire [9:0] mem_0_10_W0_addr; // @[:anonymous source@603.4]
  wire  mem_0_10_W0_clk; // @[:anonymous source@603.4]
  wire [7:0] mem_0_10_W0_data; // @[:anonymous source@603.4]
  wire  mem_0_10_W0_en; // @[:anonymous source@603.4]
  wire  mem_0_10_W0_mask; // @[:anonymous source@603.4]
  wire [9:0] mem_0_10_R0_addr; // @[:anonymous source@603.4]
  wire  mem_0_10_R0_clk; // @[:anonymous source@603.4]
  wire [7:0] mem_0_10_R0_data; // @[:anonymous source@603.4]
  wire  mem_0_10_R0_en; // @[:anonymous source@603.4]
  wire [9:0] mem_0_11_W0_addr; // @[:anonymous source@604.4]
  wire  mem_0_11_W0_clk; // @[:anonymous source@604.4]
  wire [7:0] mem_0_11_W0_data; // @[:anonymous source@604.4]
  wire  mem_0_11_W0_en; // @[:anonymous source@604.4]
  wire  mem_0_11_W0_mask; // @[:anonymous source@604.4]
  wire [9:0] mem_0_11_R0_addr; // @[:anonymous source@604.4]
  wire  mem_0_11_R0_clk; // @[:anonymous source@604.4]
  wire [7:0] mem_0_11_R0_data; // @[:anonymous source@604.4]
  wire  mem_0_11_R0_en; // @[:anonymous source@604.4]
  wire [9:0] mem_0_12_W0_addr; // @[:anonymous source@605.4]
  wire  mem_0_12_W0_clk; // @[:anonymous source@605.4]
  wire [7:0] mem_0_12_W0_data; // @[:anonymous source@605.4]
  wire  mem_0_12_W0_en; // @[:anonymous source@605.4]
  wire  mem_0_12_W0_mask; // @[:anonymous source@605.4]
  wire [9:0] mem_0_12_R0_addr; // @[:anonymous source@605.4]
  wire  mem_0_12_R0_clk; // @[:anonymous source@605.4]
  wire [7:0] mem_0_12_R0_data; // @[:anonymous source@605.4]
  wire  mem_0_12_R0_en; // @[:anonymous source@605.4]
  wire [9:0] mem_0_13_W0_addr; // @[:anonymous source@606.4]
  wire  mem_0_13_W0_clk; // @[:anonymous source@606.4]
  wire [7:0] mem_0_13_W0_data; // @[:anonymous source@606.4]
  wire  mem_0_13_W0_en; // @[:anonymous source@606.4]
  wire  mem_0_13_W0_mask; // @[:anonymous source@606.4]
  wire [9:0] mem_0_13_R0_addr; // @[:anonymous source@606.4]
  wire  mem_0_13_R0_clk; // @[:anonymous source@606.4]
  wire [7:0] mem_0_13_R0_data; // @[:anonymous source@606.4]
  wire  mem_0_13_R0_en; // @[:anonymous source@606.4]
  wire [9:0] mem_0_14_W0_addr; // @[:anonymous source@607.4]
  wire  mem_0_14_W0_clk; // @[:anonymous source@607.4]
  wire [7:0] mem_0_14_W0_data; // @[:anonymous source@607.4]
  wire  mem_0_14_W0_en; // @[:anonymous source@607.4]
  wire  mem_0_14_W0_mask; // @[:anonymous source@607.4]
  wire [9:0] mem_0_14_R0_addr; // @[:anonymous source@607.4]
  wire  mem_0_14_R0_clk; // @[:anonymous source@607.4]
  wire [7:0] mem_0_14_R0_data; // @[:anonymous source@607.4]
  wire  mem_0_14_R0_en; // @[:anonymous source@607.4]
  wire [9:0] mem_0_15_W0_addr; // @[:anonymous source@608.4]
  wire  mem_0_15_W0_clk; // @[:anonymous source@608.4]
  wire [7:0] mem_0_15_W0_data; // @[:anonymous source@608.4]
  wire  mem_0_15_W0_en; // @[:anonymous source@608.4]
  wire  mem_0_15_W0_mask; // @[:anonymous source@608.4]
  wire [9:0] mem_0_15_R0_addr; // @[:anonymous source@608.4]
  wire  mem_0_15_R0_clk; // @[:anonymous source@608.4]
  wire [7:0] mem_0_15_R0_data; // @[:anonymous source@608.4]
  wire  mem_0_15_R0_en; // @[:anonymous source@608.4]
  wire [9:0] mem_0_16_W0_addr; // @[:anonymous source@609.4]
  wire  mem_0_16_W0_clk; // @[:anonymous source@609.4]
  wire [7:0] mem_0_16_W0_data; // @[:anonymous source@609.4]
  wire  mem_0_16_W0_en; // @[:anonymous source@609.4]
  wire  mem_0_16_W0_mask; // @[:anonymous source@609.4]
  wire [9:0] mem_0_16_R0_addr; // @[:anonymous source@609.4]
  wire  mem_0_16_R0_clk; // @[:anonymous source@609.4]
  wire [7:0] mem_0_16_R0_data; // @[:anonymous source@609.4]
  wire  mem_0_16_R0_en; // @[:anonymous source@609.4]
  wire [9:0] mem_0_17_W0_addr; // @[:anonymous source@610.4]
  wire  mem_0_17_W0_clk; // @[:anonymous source@610.4]
  wire [7:0] mem_0_17_W0_data; // @[:anonymous source@610.4]
  wire  mem_0_17_W0_en; // @[:anonymous source@610.4]
  wire  mem_0_17_W0_mask; // @[:anonymous source@610.4]
  wire [9:0] mem_0_17_R0_addr; // @[:anonymous source@610.4]
  wire  mem_0_17_R0_clk; // @[:anonymous source@610.4]
  wire [7:0] mem_0_17_R0_data; // @[:anonymous source@610.4]
  wire  mem_0_17_R0_en; // @[:anonymous source@610.4]
  wire [9:0] mem_0_18_W0_addr; // @[:anonymous source@611.4]
  wire  mem_0_18_W0_clk; // @[:anonymous source@611.4]
  wire [7:0] mem_0_18_W0_data; // @[:anonymous source@611.4]
  wire  mem_0_18_W0_en; // @[:anonymous source@611.4]
  wire  mem_0_18_W0_mask; // @[:anonymous source@611.4]
  wire [9:0] mem_0_18_R0_addr; // @[:anonymous source@611.4]
  wire  mem_0_18_R0_clk; // @[:anonymous source@611.4]
  wire [7:0] mem_0_18_R0_data; // @[:anonymous source@611.4]
  wire  mem_0_18_R0_en; // @[:anonymous source@611.4]
  wire [9:0] mem_0_19_W0_addr; // @[:anonymous source@612.4]
  wire  mem_0_19_W0_clk; // @[:anonymous source@612.4]
  wire [7:0] mem_0_19_W0_data; // @[:anonymous source@612.4]
  wire  mem_0_19_W0_en; // @[:anonymous source@612.4]
  wire  mem_0_19_W0_mask; // @[:anonymous source@612.4]
  wire [9:0] mem_0_19_R0_addr; // @[:anonymous source@612.4]
  wire  mem_0_19_R0_clk; // @[:anonymous source@612.4]
  wire [7:0] mem_0_19_R0_data; // @[:anonymous source@612.4]
  wire  mem_0_19_R0_en; // @[:anonymous source@612.4]
  wire [9:0] mem_0_20_W0_addr; // @[:anonymous source@613.4]
  wire  mem_0_20_W0_clk; // @[:anonymous source@613.4]
  wire [7:0] mem_0_20_W0_data; // @[:anonymous source@613.4]
  wire  mem_0_20_W0_en; // @[:anonymous source@613.4]
  wire  mem_0_20_W0_mask; // @[:anonymous source@613.4]
  wire [9:0] mem_0_20_R0_addr; // @[:anonymous source@613.4]
  wire  mem_0_20_R0_clk; // @[:anonymous source@613.4]
  wire [7:0] mem_0_20_R0_data; // @[:anonymous source@613.4]
  wire  mem_0_20_R0_en; // @[:anonymous source@613.4]
  wire [9:0] mem_0_21_W0_addr; // @[:anonymous source@614.4]
  wire  mem_0_21_W0_clk; // @[:anonymous source@614.4]
  wire [7:0] mem_0_21_W0_data; // @[:anonymous source@614.4]
  wire  mem_0_21_W0_en; // @[:anonymous source@614.4]
  wire  mem_0_21_W0_mask; // @[:anonymous source@614.4]
  wire [9:0] mem_0_21_R0_addr; // @[:anonymous source@614.4]
  wire  mem_0_21_R0_clk; // @[:anonymous source@614.4]
  wire [7:0] mem_0_21_R0_data; // @[:anonymous source@614.4]
  wire  mem_0_21_R0_en; // @[:anonymous source@614.4]
  wire [9:0] mem_0_22_W0_addr; // @[:anonymous source@615.4]
  wire  mem_0_22_W0_clk; // @[:anonymous source@615.4]
  wire [7:0] mem_0_22_W0_data; // @[:anonymous source@615.4]
  wire  mem_0_22_W0_en; // @[:anonymous source@615.4]
  wire  mem_0_22_W0_mask; // @[:anonymous source@615.4]
  wire [9:0] mem_0_22_R0_addr; // @[:anonymous source@615.4]
  wire  mem_0_22_R0_clk; // @[:anonymous source@615.4]
  wire [7:0] mem_0_22_R0_data; // @[:anonymous source@615.4]
  wire  mem_0_22_R0_en; // @[:anonymous source@615.4]
  wire [9:0] mem_0_23_W0_addr; // @[:anonymous source@616.4]
  wire  mem_0_23_W0_clk; // @[:anonymous source@616.4]
  wire [7:0] mem_0_23_W0_data; // @[:anonymous source@616.4]
  wire  mem_0_23_W0_en; // @[:anonymous source@616.4]
  wire  mem_0_23_W0_mask; // @[:anonymous source@616.4]
  wire [9:0] mem_0_23_R0_addr; // @[:anonymous source@616.4]
  wire  mem_0_23_R0_clk; // @[:anonymous source@616.4]
  wire [7:0] mem_0_23_R0_data; // @[:anonymous source@616.4]
  wire  mem_0_23_R0_en; // @[:anonymous source@616.4]
  wire [9:0] mem_0_24_W0_addr; // @[:anonymous source@617.4]
  wire  mem_0_24_W0_clk; // @[:anonymous source@617.4]
  wire [7:0] mem_0_24_W0_data; // @[:anonymous source@617.4]
  wire  mem_0_24_W0_en; // @[:anonymous source@617.4]
  wire  mem_0_24_W0_mask; // @[:anonymous source@617.4]
  wire [9:0] mem_0_24_R0_addr; // @[:anonymous source@617.4]
  wire  mem_0_24_R0_clk; // @[:anonymous source@617.4]
  wire [7:0] mem_0_24_R0_data; // @[:anonymous source@617.4]
  wire  mem_0_24_R0_en; // @[:anonymous source@617.4]
  wire [9:0] mem_0_25_W0_addr; // @[:anonymous source@618.4]
  wire  mem_0_25_W0_clk; // @[:anonymous source@618.4]
  wire [7:0] mem_0_25_W0_data; // @[:anonymous source@618.4]
  wire  mem_0_25_W0_en; // @[:anonymous source@618.4]
  wire  mem_0_25_W0_mask; // @[:anonymous source@618.4]
  wire [9:0] mem_0_25_R0_addr; // @[:anonymous source@618.4]
  wire  mem_0_25_R0_clk; // @[:anonymous source@618.4]
  wire [7:0] mem_0_25_R0_data; // @[:anonymous source@618.4]
  wire  mem_0_25_R0_en; // @[:anonymous source@618.4]
  wire [9:0] mem_0_26_W0_addr; // @[:anonymous source@619.4]
  wire  mem_0_26_W0_clk; // @[:anonymous source@619.4]
  wire [7:0] mem_0_26_W0_data; // @[:anonymous source@619.4]
  wire  mem_0_26_W0_en; // @[:anonymous source@619.4]
  wire  mem_0_26_W0_mask; // @[:anonymous source@619.4]
  wire [9:0] mem_0_26_R0_addr; // @[:anonymous source@619.4]
  wire  mem_0_26_R0_clk; // @[:anonymous source@619.4]
  wire [7:0] mem_0_26_R0_data; // @[:anonymous source@619.4]
  wire  mem_0_26_R0_en; // @[:anonymous source@619.4]
  wire [9:0] mem_0_27_W0_addr; // @[:anonymous source@620.4]
  wire  mem_0_27_W0_clk; // @[:anonymous source@620.4]
  wire [7:0] mem_0_27_W0_data; // @[:anonymous source@620.4]
  wire  mem_0_27_W0_en; // @[:anonymous source@620.4]
  wire  mem_0_27_W0_mask; // @[:anonymous source@620.4]
  wire [9:0] mem_0_27_R0_addr; // @[:anonymous source@620.4]
  wire  mem_0_27_R0_clk; // @[:anonymous source@620.4]
  wire [7:0] mem_0_27_R0_data; // @[:anonymous source@620.4]
  wire  mem_0_27_R0_en; // @[:anonymous source@620.4]
  wire [9:0] mem_0_28_W0_addr; // @[:anonymous source@621.4]
  wire  mem_0_28_W0_clk; // @[:anonymous source@621.4]
  wire [7:0] mem_0_28_W0_data; // @[:anonymous source@621.4]
  wire  mem_0_28_W0_en; // @[:anonymous source@621.4]
  wire  mem_0_28_W0_mask; // @[:anonymous source@621.4]
  wire [9:0] mem_0_28_R0_addr; // @[:anonymous source@621.4]
  wire  mem_0_28_R0_clk; // @[:anonymous source@621.4]
  wire [7:0] mem_0_28_R0_data; // @[:anonymous source@621.4]
  wire  mem_0_28_R0_en; // @[:anonymous source@621.4]
  wire [9:0] mem_0_29_W0_addr; // @[:anonymous source@622.4]
  wire  mem_0_29_W0_clk; // @[:anonymous source@622.4]
  wire [7:0] mem_0_29_W0_data; // @[:anonymous source@622.4]
  wire  mem_0_29_W0_en; // @[:anonymous source@622.4]
  wire  mem_0_29_W0_mask; // @[:anonymous source@622.4]
  wire [9:0] mem_0_29_R0_addr; // @[:anonymous source@622.4]
  wire  mem_0_29_R0_clk; // @[:anonymous source@622.4]
  wire [7:0] mem_0_29_R0_data; // @[:anonymous source@622.4]
  wire  mem_0_29_R0_en; // @[:anonymous source@622.4]
  wire [9:0] mem_0_30_W0_addr; // @[:anonymous source@623.4]
  wire  mem_0_30_W0_clk; // @[:anonymous source@623.4]
  wire [7:0] mem_0_30_W0_data; // @[:anonymous source@623.4]
  wire  mem_0_30_W0_en; // @[:anonymous source@623.4]
  wire  mem_0_30_W0_mask; // @[:anonymous source@623.4]
  wire [9:0] mem_0_30_R0_addr; // @[:anonymous source@623.4]
  wire  mem_0_30_R0_clk; // @[:anonymous source@623.4]
  wire [7:0] mem_0_30_R0_data; // @[:anonymous source@623.4]
  wire  mem_0_30_R0_en; // @[:anonymous source@623.4]
  wire [9:0] mem_0_31_W0_addr; // @[:anonymous source@624.4]
  wire  mem_0_31_W0_clk; // @[:anonymous source@624.4]
  wire [7:0] mem_0_31_W0_data; // @[:anonymous source@624.4]
  wire  mem_0_31_W0_en; // @[:anonymous source@624.4]
  wire  mem_0_31_W0_mask; // @[:anonymous source@624.4]
  wire [9:0] mem_0_31_R0_addr; // @[:anonymous source@624.4]
  wire  mem_0_31_R0_clk; // @[:anonymous source@624.4]
  wire [7:0] mem_0_31_R0_data; // @[:anonymous source@624.4]
  wire  mem_0_31_R0_en; // @[:anonymous source@624.4]
  wire [9:0] mem_0_32_W0_addr; // @[:anonymous source@625.4]
  wire  mem_0_32_W0_clk; // @[:anonymous source@625.4]
  wire [7:0] mem_0_32_W0_data; // @[:anonymous source@625.4]
  wire  mem_0_32_W0_en; // @[:anonymous source@625.4]
  wire  mem_0_32_W0_mask; // @[:anonymous source@625.4]
  wire [9:0] mem_0_32_R0_addr; // @[:anonymous source@625.4]
  wire  mem_0_32_R0_clk; // @[:anonymous source@625.4]
  wire [7:0] mem_0_32_R0_data; // @[:anonymous source@625.4]
  wire  mem_0_32_R0_en; // @[:anonymous source@625.4]
  wire [9:0] mem_0_33_W0_addr; // @[:anonymous source@626.4]
  wire  mem_0_33_W0_clk; // @[:anonymous source@626.4]
  wire [7:0] mem_0_33_W0_data; // @[:anonymous source@626.4]
  wire  mem_0_33_W0_en; // @[:anonymous source@626.4]
  wire  mem_0_33_W0_mask; // @[:anonymous source@626.4]
  wire [9:0] mem_0_33_R0_addr; // @[:anonymous source@626.4]
  wire  mem_0_33_R0_clk; // @[:anonymous source@626.4]
  wire [7:0] mem_0_33_R0_data; // @[:anonymous source@626.4]
  wire  mem_0_33_R0_en; // @[:anonymous source@626.4]
  wire [9:0] mem_0_34_W0_addr; // @[:anonymous source@627.4]
  wire  mem_0_34_W0_clk; // @[:anonymous source@627.4]
  wire [7:0] mem_0_34_W0_data; // @[:anonymous source@627.4]
  wire  mem_0_34_W0_en; // @[:anonymous source@627.4]
  wire  mem_0_34_W0_mask; // @[:anonymous source@627.4]
  wire [9:0] mem_0_34_R0_addr; // @[:anonymous source@627.4]
  wire  mem_0_34_R0_clk; // @[:anonymous source@627.4]
  wire [7:0] mem_0_34_R0_data; // @[:anonymous source@627.4]
  wire  mem_0_34_R0_en; // @[:anonymous source@627.4]
  wire [9:0] mem_0_35_W0_addr; // @[:anonymous source@628.4]
  wire  mem_0_35_W0_clk; // @[:anonymous source@628.4]
  wire [7:0] mem_0_35_W0_data; // @[:anonymous source@628.4]
  wire  mem_0_35_W0_en; // @[:anonymous source@628.4]
  wire  mem_0_35_W0_mask; // @[:anonymous source@628.4]
  wire [9:0] mem_0_35_R0_addr; // @[:anonymous source@628.4]
  wire  mem_0_35_R0_clk; // @[:anonymous source@628.4]
  wire [7:0] mem_0_35_R0_data; // @[:anonymous source@628.4]
  wire  mem_0_35_R0_en; // @[:anonymous source@628.4]
  wire [9:0] mem_0_36_W0_addr; // @[:anonymous source@629.4]
  wire  mem_0_36_W0_clk; // @[:anonymous source@629.4]
  wire [7:0] mem_0_36_W0_data; // @[:anonymous source@629.4]
  wire  mem_0_36_W0_en; // @[:anonymous source@629.4]
  wire  mem_0_36_W0_mask; // @[:anonymous source@629.4]
  wire [9:0] mem_0_36_R0_addr; // @[:anonymous source@629.4]
  wire  mem_0_36_R0_clk; // @[:anonymous source@629.4]
  wire [7:0] mem_0_36_R0_data; // @[:anonymous source@629.4]
  wire  mem_0_36_R0_en; // @[:anonymous source@629.4]
  wire [9:0] mem_0_37_W0_addr; // @[:anonymous source@630.4]
  wire  mem_0_37_W0_clk; // @[:anonymous source@630.4]
  wire [7:0] mem_0_37_W0_data; // @[:anonymous source@630.4]
  wire  mem_0_37_W0_en; // @[:anonymous source@630.4]
  wire  mem_0_37_W0_mask; // @[:anonymous source@630.4]
  wire [9:0] mem_0_37_R0_addr; // @[:anonymous source@630.4]
  wire  mem_0_37_R0_clk; // @[:anonymous source@630.4]
  wire [7:0] mem_0_37_R0_data; // @[:anonymous source@630.4]
  wire  mem_0_37_R0_en; // @[:anonymous source@630.4]
  wire [9:0] mem_0_38_W0_addr; // @[:anonymous source@631.4]
  wire  mem_0_38_W0_clk; // @[:anonymous source@631.4]
  wire [7:0] mem_0_38_W0_data; // @[:anonymous source@631.4]
  wire  mem_0_38_W0_en; // @[:anonymous source@631.4]
  wire  mem_0_38_W0_mask; // @[:anonymous source@631.4]
  wire [9:0] mem_0_38_R0_addr; // @[:anonymous source@631.4]
  wire  mem_0_38_R0_clk; // @[:anonymous source@631.4]
  wire [7:0] mem_0_38_R0_data; // @[:anonymous source@631.4]
  wire  mem_0_38_R0_en; // @[:anonymous source@631.4]
  wire [9:0] mem_0_39_W0_addr; // @[:anonymous source@632.4]
  wire  mem_0_39_W0_clk; // @[:anonymous source@632.4]
  wire [7:0] mem_0_39_W0_data; // @[:anonymous source@632.4]
  wire  mem_0_39_W0_en; // @[:anonymous source@632.4]
  wire  mem_0_39_W0_mask; // @[:anonymous source@632.4]
  wire [9:0] mem_0_39_R0_addr; // @[:anonymous source@632.4]
  wire  mem_0_39_R0_clk; // @[:anonymous source@632.4]
  wire [7:0] mem_0_39_R0_data; // @[:anonymous source@632.4]
  wire  mem_0_39_R0_en; // @[:anonymous source@632.4]
  wire [9:0] mem_0_40_W0_addr; // @[:anonymous source@633.4]
  wire  mem_0_40_W0_clk; // @[:anonymous source@633.4]
  wire [7:0] mem_0_40_W0_data; // @[:anonymous source@633.4]
  wire  mem_0_40_W0_en; // @[:anonymous source@633.4]
  wire  mem_0_40_W0_mask; // @[:anonymous source@633.4]
  wire [9:0] mem_0_40_R0_addr; // @[:anonymous source@633.4]
  wire  mem_0_40_R0_clk; // @[:anonymous source@633.4]
  wire [7:0] mem_0_40_R0_data; // @[:anonymous source@633.4]
  wire  mem_0_40_R0_en; // @[:anonymous source@633.4]
  wire [9:0] mem_0_41_W0_addr; // @[:anonymous source@634.4]
  wire  mem_0_41_W0_clk; // @[:anonymous source@634.4]
  wire [7:0] mem_0_41_W0_data; // @[:anonymous source@634.4]
  wire  mem_0_41_W0_en; // @[:anonymous source@634.4]
  wire  mem_0_41_W0_mask; // @[:anonymous source@634.4]
  wire [9:0] mem_0_41_R0_addr; // @[:anonymous source@634.4]
  wire  mem_0_41_R0_clk; // @[:anonymous source@634.4]
  wire [7:0] mem_0_41_R0_data; // @[:anonymous source@634.4]
  wire  mem_0_41_R0_en; // @[:anonymous source@634.4]
  wire [9:0] mem_0_42_W0_addr; // @[:anonymous source@635.4]
  wire  mem_0_42_W0_clk; // @[:anonymous source@635.4]
  wire [7:0] mem_0_42_W0_data; // @[:anonymous source@635.4]
  wire  mem_0_42_W0_en; // @[:anonymous source@635.4]
  wire  mem_0_42_W0_mask; // @[:anonymous source@635.4]
  wire [9:0] mem_0_42_R0_addr; // @[:anonymous source@635.4]
  wire  mem_0_42_R0_clk; // @[:anonymous source@635.4]
  wire [7:0] mem_0_42_R0_data; // @[:anonymous source@635.4]
  wire  mem_0_42_R0_en; // @[:anonymous source@635.4]
  wire [9:0] mem_0_43_W0_addr; // @[:anonymous source@636.4]
  wire  mem_0_43_W0_clk; // @[:anonymous source@636.4]
  wire [7:0] mem_0_43_W0_data; // @[:anonymous source@636.4]
  wire  mem_0_43_W0_en; // @[:anonymous source@636.4]
  wire  mem_0_43_W0_mask; // @[:anonymous source@636.4]
  wire [9:0] mem_0_43_R0_addr; // @[:anonymous source@636.4]
  wire  mem_0_43_R0_clk; // @[:anonymous source@636.4]
  wire [7:0] mem_0_43_R0_data; // @[:anonymous source@636.4]
  wire  mem_0_43_R0_en; // @[:anonymous source@636.4]
  wire [9:0] mem_0_44_W0_addr; // @[:anonymous source@637.4]
  wire  mem_0_44_W0_clk; // @[:anonymous source@637.4]
  wire [7:0] mem_0_44_W0_data; // @[:anonymous source@637.4]
  wire  mem_0_44_W0_en; // @[:anonymous source@637.4]
  wire  mem_0_44_W0_mask; // @[:anonymous source@637.4]
  wire [9:0] mem_0_44_R0_addr; // @[:anonymous source@637.4]
  wire  mem_0_44_R0_clk; // @[:anonymous source@637.4]
  wire [7:0] mem_0_44_R0_data; // @[:anonymous source@637.4]
  wire  mem_0_44_R0_en; // @[:anonymous source@637.4]
  wire [9:0] mem_0_45_W0_addr; // @[:anonymous source@638.4]
  wire  mem_0_45_W0_clk; // @[:anonymous source@638.4]
  wire [7:0] mem_0_45_W0_data; // @[:anonymous source@638.4]
  wire  mem_0_45_W0_en; // @[:anonymous source@638.4]
  wire  mem_0_45_W0_mask; // @[:anonymous source@638.4]
  wire [9:0] mem_0_45_R0_addr; // @[:anonymous source@638.4]
  wire  mem_0_45_R0_clk; // @[:anonymous source@638.4]
  wire [7:0] mem_0_45_R0_data; // @[:anonymous source@638.4]
  wire  mem_0_45_R0_en; // @[:anonymous source@638.4]
  wire [9:0] mem_0_46_W0_addr; // @[:anonymous source@639.4]
  wire  mem_0_46_W0_clk; // @[:anonymous source@639.4]
  wire [7:0] mem_0_46_W0_data; // @[:anonymous source@639.4]
  wire  mem_0_46_W0_en; // @[:anonymous source@639.4]
  wire  mem_0_46_W0_mask; // @[:anonymous source@639.4]
  wire [9:0] mem_0_46_R0_addr; // @[:anonymous source@639.4]
  wire  mem_0_46_R0_clk; // @[:anonymous source@639.4]
  wire [7:0] mem_0_46_R0_data; // @[:anonymous source@639.4]
  wire  mem_0_46_R0_en; // @[:anonymous source@639.4]
  wire [9:0] mem_0_47_W0_addr; // @[:anonymous source@640.4]
  wire  mem_0_47_W0_clk; // @[:anonymous source@640.4]
  wire [7:0] mem_0_47_W0_data; // @[:anonymous source@640.4]
  wire  mem_0_47_W0_en; // @[:anonymous source@640.4]
  wire  mem_0_47_W0_mask; // @[:anonymous source@640.4]
  wire [9:0] mem_0_47_R0_addr; // @[:anonymous source@640.4]
  wire  mem_0_47_R0_clk; // @[:anonymous source@640.4]
  wire [7:0] mem_0_47_R0_data; // @[:anonymous source@640.4]
  wire  mem_0_47_R0_en; // @[:anonymous source@640.4]
  wire [9:0] mem_0_48_W0_addr; // @[:anonymous source@641.4]
  wire  mem_0_48_W0_clk; // @[:anonymous source@641.4]
  wire [7:0] mem_0_48_W0_data; // @[:anonymous source@641.4]
  wire  mem_0_48_W0_en; // @[:anonymous source@641.4]
  wire  mem_0_48_W0_mask; // @[:anonymous source@641.4]
  wire [9:0] mem_0_48_R0_addr; // @[:anonymous source@641.4]
  wire  mem_0_48_R0_clk; // @[:anonymous source@641.4]
  wire [7:0] mem_0_48_R0_data; // @[:anonymous source@641.4]
  wire  mem_0_48_R0_en; // @[:anonymous source@641.4]
  wire [9:0] mem_0_49_W0_addr; // @[:anonymous source@642.4]
  wire  mem_0_49_W0_clk; // @[:anonymous source@642.4]
  wire [7:0] mem_0_49_W0_data; // @[:anonymous source@642.4]
  wire  mem_0_49_W0_en; // @[:anonymous source@642.4]
  wire  mem_0_49_W0_mask; // @[:anonymous source@642.4]
  wire [9:0] mem_0_49_R0_addr; // @[:anonymous source@642.4]
  wire  mem_0_49_R0_clk; // @[:anonymous source@642.4]
  wire [7:0] mem_0_49_R0_data; // @[:anonymous source@642.4]
  wire  mem_0_49_R0_en; // @[:anonymous source@642.4]
  wire [9:0] mem_0_50_W0_addr; // @[:anonymous source@643.4]
  wire  mem_0_50_W0_clk; // @[:anonymous source@643.4]
  wire [7:0] mem_0_50_W0_data; // @[:anonymous source@643.4]
  wire  mem_0_50_W0_en; // @[:anonymous source@643.4]
  wire  mem_0_50_W0_mask; // @[:anonymous source@643.4]
  wire [9:0] mem_0_50_R0_addr; // @[:anonymous source@643.4]
  wire  mem_0_50_R0_clk; // @[:anonymous source@643.4]
  wire [7:0] mem_0_50_R0_data; // @[:anonymous source@643.4]
  wire  mem_0_50_R0_en; // @[:anonymous source@643.4]
  wire [9:0] mem_0_51_W0_addr; // @[:anonymous source@644.4]
  wire  mem_0_51_W0_clk; // @[:anonymous source@644.4]
  wire [7:0] mem_0_51_W0_data; // @[:anonymous source@644.4]
  wire  mem_0_51_W0_en; // @[:anonymous source@644.4]
  wire  mem_0_51_W0_mask; // @[:anonymous source@644.4]
  wire [9:0] mem_0_51_R0_addr; // @[:anonymous source@644.4]
  wire  mem_0_51_R0_clk; // @[:anonymous source@644.4]
  wire [7:0] mem_0_51_R0_data; // @[:anonymous source@644.4]
  wire  mem_0_51_R0_en; // @[:anonymous source@644.4]
  wire [9:0] mem_0_52_W0_addr; // @[:anonymous source@645.4]
  wire  mem_0_52_W0_clk; // @[:anonymous source@645.4]
  wire [7:0] mem_0_52_W0_data; // @[:anonymous source@645.4]
  wire  mem_0_52_W0_en; // @[:anonymous source@645.4]
  wire  mem_0_52_W0_mask; // @[:anonymous source@645.4]
  wire [9:0] mem_0_52_R0_addr; // @[:anonymous source@645.4]
  wire  mem_0_52_R0_clk; // @[:anonymous source@645.4]
  wire [7:0] mem_0_52_R0_data; // @[:anonymous source@645.4]
  wire  mem_0_52_R0_en; // @[:anonymous source@645.4]
  wire [9:0] mem_0_53_W0_addr; // @[:anonymous source@646.4]
  wire  mem_0_53_W0_clk; // @[:anonymous source@646.4]
  wire [7:0] mem_0_53_W0_data; // @[:anonymous source@646.4]
  wire  mem_0_53_W0_en; // @[:anonymous source@646.4]
  wire  mem_0_53_W0_mask; // @[:anonymous source@646.4]
  wire [9:0] mem_0_53_R0_addr; // @[:anonymous source@646.4]
  wire  mem_0_53_R0_clk; // @[:anonymous source@646.4]
  wire [7:0] mem_0_53_R0_data; // @[:anonymous source@646.4]
  wire  mem_0_53_R0_en; // @[:anonymous source@646.4]
  wire [9:0] mem_0_54_W0_addr; // @[:anonymous source@647.4]
  wire  mem_0_54_W0_clk; // @[:anonymous source@647.4]
  wire [7:0] mem_0_54_W0_data; // @[:anonymous source@647.4]
  wire  mem_0_54_W0_en; // @[:anonymous source@647.4]
  wire  mem_0_54_W0_mask; // @[:anonymous source@647.4]
  wire [9:0] mem_0_54_R0_addr; // @[:anonymous source@647.4]
  wire  mem_0_54_R0_clk; // @[:anonymous source@647.4]
  wire [7:0] mem_0_54_R0_data; // @[:anonymous source@647.4]
  wire  mem_0_54_R0_en; // @[:anonymous source@647.4]
  wire [9:0] mem_0_55_W0_addr; // @[:anonymous source@648.4]
  wire  mem_0_55_W0_clk; // @[:anonymous source@648.4]
  wire [7:0] mem_0_55_W0_data; // @[:anonymous source@648.4]
  wire  mem_0_55_W0_en; // @[:anonymous source@648.4]
  wire  mem_0_55_W0_mask; // @[:anonymous source@648.4]
  wire [9:0] mem_0_55_R0_addr; // @[:anonymous source@648.4]
  wire  mem_0_55_R0_clk; // @[:anonymous source@648.4]
  wire [7:0] mem_0_55_R0_data; // @[:anonymous source@648.4]
  wire  mem_0_55_R0_en; // @[:anonymous source@648.4]
  wire [9:0] mem_0_56_W0_addr; // @[:anonymous source@649.4]
  wire  mem_0_56_W0_clk; // @[:anonymous source@649.4]
  wire [7:0] mem_0_56_W0_data; // @[:anonymous source@649.4]
  wire  mem_0_56_W0_en; // @[:anonymous source@649.4]
  wire  mem_0_56_W0_mask; // @[:anonymous source@649.4]
  wire [9:0] mem_0_56_R0_addr; // @[:anonymous source@649.4]
  wire  mem_0_56_R0_clk; // @[:anonymous source@649.4]
  wire [7:0] mem_0_56_R0_data; // @[:anonymous source@649.4]
  wire  mem_0_56_R0_en; // @[:anonymous source@649.4]
  wire [9:0] mem_0_57_W0_addr; // @[:anonymous source@650.4]
  wire  mem_0_57_W0_clk; // @[:anonymous source@650.4]
  wire [7:0] mem_0_57_W0_data; // @[:anonymous source@650.4]
  wire  mem_0_57_W0_en; // @[:anonymous source@650.4]
  wire  mem_0_57_W0_mask; // @[:anonymous source@650.4]
  wire [9:0] mem_0_57_R0_addr; // @[:anonymous source@650.4]
  wire  mem_0_57_R0_clk; // @[:anonymous source@650.4]
  wire [7:0] mem_0_57_R0_data; // @[:anonymous source@650.4]
  wire  mem_0_57_R0_en; // @[:anonymous source@650.4]
  wire [9:0] mem_0_58_W0_addr; // @[:anonymous source@651.4]
  wire  mem_0_58_W0_clk; // @[:anonymous source@651.4]
  wire [7:0] mem_0_58_W0_data; // @[:anonymous source@651.4]
  wire  mem_0_58_W0_en; // @[:anonymous source@651.4]
  wire  mem_0_58_W0_mask; // @[:anonymous source@651.4]
  wire [9:0] mem_0_58_R0_addr; // @[:anonymous source@651.4]
  wire  mem_0_58_R0_clk; // @[:anonymous source@651.4]
  wire [7:0] mem_0_58_R0_data; // @[:anonymous source@651.4]
  wire  mem_0_58_R0_en; // @[:anonymous source@651.4]
  wire [9:0] mem_0_59_W0_addr; // @[:anonymous source@652.4]
  wire  mem_0_59_W0_clk; // @[:anonymous source@652.4]
  wire [7:0] mem_0_59_W0_data; // @[:anonymous source@652.4]
  wire  mem_0_59_W0_en; // @[:anonymous source@652.4]
  wire  mem_0_59_W0_mask; // @[:anonymous source@652.4]
  wire [9:0] mem_0_59_R0_addr; // @[:anonymous source@652.4]
  wire  mem_0_59_R0_clk; // @[:anonymous source@652.4]
  wire [7:0] mem_0_59_R0_data; // @[:anonymous source@652.4]
  wire  mem_0_59_R0_en; // @[:anonymous source@652.4]
  wire [9:0] mem_0_60_W0_addr; // @[:anonymous source@653.4]
  wire  mem_0_60_W0_clk; // @[:anonymous source@653.4]
  wire [7:0] mem_0_60_W0_data; // @[:anonymous source@653.4]
  wire  mem_0_60_W0_en; // @[:anonymous source@653.4]
  wire  mem_0_60_W0_mask; // @[:anonymous source@653.4]
  wire [9:0] mem_0_60_R0_addr; // @[:anonymous source@653.4]
  wire  mem_0_60_R0_clk; // @[:anonymous source@653.4]
  wire [7:0] mem_0_60_R0_data; // @[:anonymous source@653.4]
  wire  mem_0_60_R0_en; // @[:anonymous source@653.4]
  wire [9:0] mem_0_61_W0_addr; // @[:anonymous source@654.4]
  wire  mem_0_61_W0_clk; // @[:anonymous source@654.4]
  wire [7:0] mem_0_61_W0_data; // @[:anonymous source@654.4]
  wire  mem_0_61_W0_en; // @[:anonymous source@654.4]
  wire  mem_0_61_W0_mask; // @[:anonymous source@654.4]
  wire [9:0] mem_0_61_R0_addr; // @[:anonymous source@654.4]
  wire  mem_0_61_R0_clk; // @[:anonymous source@654.4]
  wire [7:0] mem_0_61_R0_data; // @[:anonymous source@654.4]
  wire  mem_0_61_R0_en; // @[:anonymous source@654.4]
  wire [9:0] mem_0_62_W0_addr; // @[:anonymous source@655.4]
  wire  mem_0_62_W0_clk; // @[:anonymous source@655.4]
  wire [7:0] mem_0_62_W0_data; // @[:anonymous source@655.4]
  wire  mem_0_62_W0_en; // @[:anonymous source@655.4]
  wire  mem_0_62_W0_mask; // @[:anonymous source@655.4]
  wire [9:0] mem_0_62_R0_addr; // @[:anonymous source@655.4]
  wire  mem_0_62_R0_clk; // @[:anonymous source@655.4]
  wire [7:0] mem_0_62_R0_data; // @[:anonymous source@655.4]
  wire  mem_0_62_R0_en; // @[:anonymous source@655.4]
  wire [9:0] mem_0_63_W0_addr; // @[:anonymous source@656.4]
  wire  mem_0_63_W0_clk; // @[:anonymous source@656.4]
  wire [7:0] mem_0_63_W0_data; // @[:anonymous source@656.4]
  wire  mem_0_63_W0_en; // @[:anonymous source@656.4]
  wire  mem_0_63_W0_mask; // @[:anonymous source@656.4]
  wire [9:0] mem_0_63_R0_addr; // @[:anonymous source@656.4]
  wire  mem_0_63_R0_clk; // @[:anonymous source@656.4]
  wire [7:0] mem_0_63_R0_data; // @[:anonymous source@656.4]
  wire  mem_0_63_R0_en; // @[:anonymous source@656.4]
  wire [7:0] R0_data_0_0; // @[:anonymous source@979.4]
  wire [7:0] R0_data_0_1; // @[:anonymous source@983.4]
  wire [7:0] R0_data_0_2; // @[:anonymous source@987.4]
  wire [7:0] R0_data_0_3; // @[:anonymous source@991.4]
  wire [7:0] R0_data_0_4; // @[:anonymous source@995.4]
  wire [7:0] R0_data_0_5; // @[:anonymous source@999.4]
  wire [7:0] R0_data_0_6; // @[:anonymous source@1003.4]
  wire [7:0] R0_data_0_7; // @[:anonymous source@1007.4]
  wire [7:0] R0_data_0_8; // @[:anonymous source@1011.4]
  wire [7:0] R0_data_0_9; // @[:anonymous source@1015.4]
  wire [7:0] R0_data_0_10; // @[:anonymous source@1019.4]
  wire [7:0] R0_data_0_11; // @[:anonymous source@1023.4]
  wire [7:0] R0_data_0_12; // @[:anonymous source@1027.4]
  wire [7:0] R0_data_0_13; // @[:anonymous source@1031.4]
  wire [7:0] R0_data_0_14; // @[:anonymous source@1035.4]
  wire [7:0] R0_data_0_15; // @[:anonymous source@1039.4]
  wire [7:0] R0_data_0_16; // @[:anonymous source@1043.4]
  wire [7:0] R0_data_0_17; // @[:anonymous source@1047.4]
  wire [7:0] R0_data_0_18; // @[:anonymous source@1051.4]
  wire [7:0] R0_data_0_19; // @[:anonymous source@1055.4]
  wire [7:0] R0_data_0_20; // @[:anonymous source@1059.4]
  wire [7:0] R0_data_0_21; // @[:anonymous source@1063.4]
  wire [7:0] R0_data_0_22; // @[:anonymous source@1067.4]
  wire [7:0] R0_data_0_23; // @[:anonymous source@1071.4]
  wire [7:0] R0_data_0_24; // @[:anonymous source@1075.4]
  wire [7:0] R0_data_0_25; // @[:anonymous source@1079.4]
  wire [7:0] R0_data_0_26; // @[:anonymous source@1083.4]
  wire [7:0] R0_data_0_27; // @[:anonymous source@1087.4]
  wire [7:0] R0_data_0_28; // @[:anonymous source@1091.4]
  wire [7:0] R0_data_0_29; // @[:anonymous source@1095.4]
  wire [7:0] R0_data_0_30; // @[:anonymous source@1099.4]
  wire [7:0] R0_data_0_31; // @[:anonymous source@1103.4]
  wire [7:0] R0_data_0_32; // @[:anonymous source@1107.4]
  wire [7:0] R0_data_0_33; // @[:anonymous source@1111.4]
  wire [7:0] R0_data_0_34; // @[:anonymous source@1115.4]
  wire [7:0] R0_data_0_35; // @[:anonymous source@1119.4]
  wire [7:0] R0_data_0_36; // @[:anonymous source@1123.4]
  wire [7:0] R0_data_0_37; // @[:anonymous source@1127.4]
  wire [7:0] R0_data_0_38; // @[:anonymous source@1131.4]
  wire [7:0] R0_data_0_39; // @[:anonymous source@1135.4]
  wire [7:0] R0_data_0_40; // @[:anonymous source@1139.4]
  wire [7:0] R0_data_0_41; // @[:anonymous source@1143.4]
  wire [7:0] R0_data_0_42; // @[:anonymous source@1147.4]
  wire [7:0] R0_data_0_43; // @[:anonymous source@1151.4]
  wire [7:0] R0_data_0_44; // @[:anonymous source@1155.4]
  wire [7:0] R0_data_0_45; // @[:anonymous source@1159.4]
  wire [7:0] R0_data_0_46; // @[:anonymous source@1163.4]
  wire [7:0] R0_data_0_47; // @[:anonymous source@1167.4]
  wire [7:0] R0_data_0_48; // @[:anonymous source@1171.4]
  wire [7:0] R0_data_0_49; // @[:anonymous source@1175.4]
  wire [7:0] R0_data_0_50; // @[:anonymous source@1179.4]
  wire [7:0] R0_data_0_51; // @[:anonymous source@1183.4]
  wire [7:0] R0_data_0_52; // @[:anonymous source@1187.4]
  wire [7:0] R0_data_0_53; // @[:anonymous source@1191.4]
  wire [7:0] R0_data_0_54; // @[:anonymous source@1195.4]
  wire [7:0] R0_data_0_55; // @[:anonymous source@1199.4]
  wire [7:0] R0_data_0_56; // @[:anonymous source@1203.4]
  wire [7:0] R0_data_0_57; // @[:anonymous source@1207.4]
  wire [7:0] R0_data_0_58; // @[:anonymous source@1211.4]
  wire [7:0] R0_data_0_59; // @[:anonymous source@1215.4]
  wire [7:0] R0_data_0_60; // @[:anonymous source@1219.4]
  wire [7:0] R0_data_0_61; // @[:anonymous source@1223.4]
  wire [7:0] R0_data_0_62; // @[:anonymous source@1227.4]
  wire [7:0] R0_data_0_63; // @[:anonymous source@1231.4]
  wire [15:0] _GEN_0; // @[:anonymous source@1233.4]
  wire [23:0] _GEN_1; // @[:anonymous source@1233.4]
  wire [31:0] _GEN_2; // @[:anonymous source@1233.4]
  wire [39:0] _GEN_3; // @[:anonymous source@1233.4]
  wire [47:0] _GEN_4; // @[:anonymous source@1233.4]
  wire [55:0] _GEN_5; // @[:anonymous source@1233.4]
  wire [63:0] _GEN_6; // @[:anonymous source@1233.4]
  wire [71:0] _GEN_7; // @[:anonymous source@1233.4]
  wire [79:0] _GEN_8; // @[:anonymous source@1233.4]
  wire [87:0] _GEN_9; // @[:anonymous source@1233.4]
  wire [95:0] _GEN_10; // @[:anonymous source@1233.4]
  wire [103:0] _GEN_11; // @[:anonymous source@1233.4]
  wire [111:0] _GEN_12; // @[:anonymous source@1233.4]
  wire [119:0] _GEN_13; // @[:anonymous source@1233.4]
  wire [127:0] _GEN_14; // @[:anonymous source@1233.4]
  wire [135:0] _GEN_15; // @[:anonymous source@1233.4]
  wire [143:0] _GEN_16; // @[:anonymous source@1233.4]
  wire [151:0] _GEN_17; // @[:anonymous source@1233.4]
  wire [159:0] _GEN_18; // @[:anonymous source@1233.4]
  wire [167:0] _GEN_19; // @[:anonymous source@1233.4]
  wire [175:0] _GEN_20; // @[:anonymous source@1233.4]
  wire [183:0] _GEN_21; // @[:anonymous source@1233.4]
  wire [191:0] _GEN_22; // @[:anonymous source@1233.4]
  wire [199:0] _GEN_23; // @[:anonymous source@1233.4]
  wire [207:0] _GEN_24; // @[:anonymous source@1233.4]
  wire [215:0] _GEN_25; // @[:anonymous source@1233.4]
  wire [223:0] _GEN_26; // @[:anonymous source@1233.4]
  wire [231:0] _GEN_27; // @[:anonymous source@1233.4]
  wire [239:0] _GEN_28; // @[:anonymous source@1233.4]
  wire [247:0] _GEN_29; // @[:anonymous source@1233.4]
  wire [255:0] _GEN_30; // @[:anonymous source@1233.4]
  wire [263:0] _GEN_31; // @[:anonymous source@1233.4]
  wire [271:0] _GEN_32; // @[:anonymous source@1233.4]
  wire [279:0] _GEN_33; // @[:anonymous source@1233.4]
  wire [287:0] _GEN_34; // @[:anonymous source@1233.4]
  wire [295:0] _GEN_35; // @[:anonymous source@1233.4]
  wire [303:0] _GEN_36; // @[:anonymous source@1233.4]
  wire [311:0] _GEN_37; // @[:anonymous source@1233.4]
  wire [319:0] _GEN_38; // @[:anonymous source@1233.4]
  wire [327:0] _GEN_39; // @[:anonymous source@1233.4]
  wire [335:0] _GEN_40; // @[:anonymous source@1233.4]
  wire [343:0] _GEN_41; // @[:anonymous source@1233.4]
  wire [351:0] _GEN_42; // @[:anonymous source@1233.4]
  wire [359:0] _GEN_43; // @[:anonymous source@1233.4]
  wire [367:0] _GEN_44; // @[:anonymous source@1233.4]
  wire [375:0] _GEN_45; // @[:anonymous source@1233.4]
  wire [383:0] _GEN_46; // @[:anonymous source@1233.4]
  wire [391:0] _GEN_47; // @[:anonymous source@1233.4]
  wire [399:0] _GEN_48; // @[:anonymous source@1233.4]
  wire [407:0] _GEN_49; // @[:anonymous source@1233.4]
  wire [415:0] _GEN_50; // @[:anonymous source@1233.4]
  wire [423:0] _GEN_51; // @[:anonymous source@1233.4]
  wire [431:0] _GEN_52; // @[:anonymous source@1233.4]
  wire [439:0] _GEN_53; // @[:anonymous source@1233.4]
  wire [447:0] _GEN_54; // @[:anonymous source@1233.4]
  wire [455:0] _GEN_55; // @[:anonymous source@1233.4]
  wire [463:0] _GEN_56; // @[:anonymous source@1233.4]
  wire [471:0] _GEN_57; // @[:anonymous source@1233.4]
  wire [479:0] _GEN_58; // @[:anonymous source@1233.4]
  wire [487:0] _GEN_59; // @[:anonymous source@1233.4]
  wire [495:0] _GEN_60; // @[:anonymous source@1233.4]
  wire [503:0] _GEN_61; // @[:anonymous source@1233.4]
  wire [511:0] R0_data_0; // @[:anonymous source@1233.4]
  wire [15:0] _GEN_62; // @[:anonymous source@1234.4]
  wire [23:0] _GEN_63; // @[:anonymous source@1234.4]
  wire [31:0] _GEN_64; // @[:anonymous source@1234.4]
  wire [39:0] _GEN_65; // @[:anonymous source@1234.4]
  wire [47:0] _GEN_66; // @[:anonymous source@1234.4]
  wire [55:0] _GEN_67; // @[:anonymous source@1234.4]
  wire [63:0] _GEN_68; // @[:anonymous source@1234.4]
  wire [71:0] _GEN_69; // @[:anonymous source@1234.4]
  wire [79:0] _GEN_70; // @[:anonymous source@1234.4]
  wire [87:0] _GEN_71; // @[:anonymous source@1234.4]
  wire [95:0] _GEN_72; // @[:anonymous source@1234.4]
  wire [103:0] _GEN_73; // @[:anonymous source@1234.4]
  wire [111:0] _GEN_74; // @[:anonymous source@1234.4]
  wire [119:0] _GEN_75; // @[:anonymous source@1234.4]
  wire [127:0] _GEN_76; // @[:anonymous source@1234.4]
  wire [135:0] _GEN_77; // @[:anonymous source@1234.4]
  wire [143:0] _GEN_78; // @[:anonymous source@1234.4]
  wire [151:0] _GEN_79; // @[:anonymous source@1234.4]
  wire [159:0] _GEN_80; // @[:anonymous source@1234.4]
  wire [167:0] _GEN_81; // @[:anonymous source@1234.4]
  wire [175:0] _GEN_82; // @[:anonymous source@1234.4]
  wire [183:0] _GEN_83; // @[:anonymous source@1234.4]
  wire [191:0] _GEN_84; // @[:anonymous source@1234.4]
  wire [199:0] _GEN_85; // @[:anonymous source@1234.4]
  wire [207:0] _GEN_86; // @[:anonymous source@1234.4]
  wire [215:0] _GEN_87; // @[:anonymous source@1234.4]
  wire [223:0] _GEN_88; // @[:anonymous source@1234.4]
  wire [231:0] _GEN_89; // @[:anonymous source@1234.4]
  wire [239:0] _GEN_90; // @[:anonymous source@1234.4]
  wire [247:0] _GEN_91; // @[:anonymous source@1234.4]
  wire [255:0] _GEN_92; // @[:anonymous source@1234.4]
  wire [263:0] _GEN_93; // @[:anonymous source@1234.4]
  wire [271:0] _GEN_94; // @[:anonymous source@1234.4]
  wire [279:0] _GEN_95; // @[:anonymous source@1234.4]
  wire [287:0] _GEN_96; // @[:anonymous source@1234.4]
  wire [295:0] _GEN_97; // @[:anonymous source@1234.4]
  wire [303:0] _GEN_98; // @[:anonymous source@1234.4]
  wire [311:0] _GEN_99; // @[:anonymous source@1234.4]
  wire [319:0] _GEN_100; // @[:anonymous source@1234.4]
  wire [327:0] _GEN_101; // @[:anonymous source@1234.4]
  wire [335:0] _GEN_102; // @[:anonymous source@1234.4]
  wire [343:0] _GEN_103; // @[:anonymous source@1234.4]
  wire [351:0] _GEN_104; // @[:anonymous source@1234.4]
  wire [359:0] _GEN_105; // @[:anonymous source@1234.4]
  wire [367:0] _GEN_106; // @[:anonymous source@1234.4]
  wire [375:0] _GEN_107; // @[:anonymous source@1234.4]
  wire [383:0] _GEN_108; // @[:anonymous source@1234.4]
  wire [391:0] _GEN_109; // @[:anonymous source@1234.4]
  wire [399:0] _GEN_110; // @[:anonymous source@1234.4]
  wire [407:0] _GEN_111; // @[:anonymous source@1234.4]
  wire [415:0] _GEN_112; // @[:anonymous source@1234.4]
  wire [423:0] _GEN_113; // @[:anonymous source@1234.4]
  wire [431:0] _GEN_114; // @[:anonymous source@1234.4]
  wire [439:0] _GEN_115; // @[:anonymous source@1234.4]
  wire [447:0] _GEN_116; // @[:anonymous source@1234.4]
  wire [455:0] _GEN_117; // @[:anonymous source@1234.4]
  wire [463:0] _GEN_118; // @[:anonymous source@1234.4]
  wire [471:0] _GEN_119; // @[:anonymous source@1234.4]
  wire [479:0] _GEN_120; // @[:anonymous source@1234.4]
  wire [487:0] _GEN_121; // @[:anonymous source@1234.4]
  wire [495:0] _GEN_122; // @[:anonymous source@1234.4]
  wire [503:0] _GEN_123; // @[:anonymous source@1234.4]
  split_mem_0_ext mem_0_0 ( // @[:anonymous source@593.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_mem_0_ext mem_0_1 ( // @[:anonymous source@594.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_mem_0_ext mem_0_2 ( // @[:anonymous source@595.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_mem_0_ext mem_0_3 ( // @[:anonymous source@596.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  split_mem_0_ext mem_0_4 ( // @[:anonymous source@597.4]
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask),
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en)
  );
  split_mem_0_ext mem_0_5 ( // @[:anonymous source@598.4]
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask),
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en)
  );
  split_mem_0_ext mem_0_6 ( // @[:anonymous source@599.4]
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask),
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en)
  );
  split_mem_0_ext mem_0_7 ( // @[:anonymous source@600.4]
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask),
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en)
  );
  split_mem_0_ext mem_0_8 ( // @[:anonymous source@601.4]
    .W0_addr(mem_0_8_W0_addr),
    .W0_clk(mem_0_8_W0_clk),
    .W0_data(mem_0_8_W0_data),
    .W0_en(mem_0_8_W0_en),
    .W0_mask(mem_0_8_W0_mask),
    .R0_addr(mem_0_8_R0_addr),
    .R0_clk(mem_0_8_R0_clk),
    .R0_data(mem_0_8_R0_data),
    .R0_en(mem_0_8_R0_en)
  );
  split_mem_0_ext mem_0_9 ( // @[:anonymous source@602.4]
    .W0_addr(mem_0_9_W0_addr),
    .W0_clk(mem_0_9_W0_clk),
    .W0_data(mem_0_9_W0_data),
    .W0_en(mem_0_9_W0_en),
    .W0_mask(mem_0_9_W0_mask),
    .R0_addr(mem_0_9_R0_addr),
    .R0_clk(mem_0_9_R0_clk),
    .R0_data(mem_0_9_R0_data),
    .R0_en(mem_0_9_R0_en)
  );
  split_mem_0_ext mem_0_10 ( // @[:anonymous source@603.4]
    .W0_addr(mem_0_10_W0_addr),
    .W0_clk(mem_0_10_W0_clk),
    .W0_data(mem_0_10_W0_data),
    .W0_en(mem_0_10_W0_en),
    .W0_mask(mem_0_10_W0_mask),
    .R0_addr(mem_0_10_R0_addr),
    .R0_clk(mem_0_10_R0_clk),
    .R0_data(mem_0_10_R0_data),
    .R0_en(mem_0_10_R0_en)
  );
  split_mem_0_ext mem_0_11 ( // @[:anonymous source@604.4]
    .W0_addr(mem_0_11_W0_addr),
    .W0_clk(mem_0_11_W0_clk),
    .W0_data(mem_0_11_W0_data),
    .W0_en(mem_0_11_W0_en),
    .W0_mask(mem_0_11_W0_mask),
    .R0_addr(mem_0_11_R0_addr),
    .R0_clk(mem_0_11_R0_clk),
    .R0_data(mem_0_11_R0_data),
    .R0_en(mem_0_11_R0_en)
  );
  split_mem_0_ext mem_0_12 ( // @[:anonymous source@605.4]
    .W0_addr(mem_0_12_W0_addr),
    .W0_clk(mem_0_12_W0_clk),
    .W0_data(mem_0_12_W0_data),
    .W0_en(mem_0_12_W0_en),
    .W0_mask(mem_0_12_W0_mask),
    .R0_addr(mem_0_12_R0_addr),
    .R0_clk(mem_0_12_R0_clk),
    .R0_data(mem_0_12_R0_data),
    .R0_en(mem_0_12_R0_en)
  );
  split_mem_0_ext mem_0_13 ( // @[:anonymous source@606.4]
    .W0_addr(mem_0_13_W0_addr),
    .W0_clk(mem_0_13_W0_clk),
    .W0_data(mem_0_13_W0_data),
    .W0_en(mem_0_13_W0_en),
    .W0_mask(mem_0_13_W0_mask),
    .R0_addr(mem_0_13_R0_addr),
    .R0_clk(mem_0_13_R0_clk),
    .R0_data(mem_0_13_R0_data),
    .R0_en(mem_0_13_R0_en)
  );
  split_mem_0_ext mem_0_14 ( // @[:anonymous source@607.4]
    .W0_addr(mem_0_14_W0_addr),
    .W0_clk(mem_0_14_W0_clk),
    .W0_data(mem_0_14_W0_data),
    .W0_en(mem_0_14_W0_en),
    .W0_mask(mem_0_14_W0_mask),
    .R0_addr(mem_0_14_R0_addr),
    .R0_clk(mem_0_14_R0_clk),
    .R0_data(mem_0_14_R0_data),
    .R0_en(mem_0_14_R0_en)
  );
  split_mem_0_ext mem_0_15 ( // @[:anonymous source@608.4]
    .W0_addr(mem_0_15_W0_addr),
    .W0_clk(mem_0_15_W0_clk),
    .W0_data(mem_0_15_W0_data),
    .W0_en(mem_0_15_W0_en),
    .W0_mask(mem_0_15_W0_mask),
    .R0_addr(mem_0_15_R0_addr),
    .R0_clk(mem_0_15_R0_clk),
    .R0_data(mem_0_15_R0_data),
    .R0_en(mem_0_15_R0_en)
  );
  split_mem_0_ext mem_0_16 ( // @[:anonymous source@609.4]
    .W0_addr(mem_0_16_W0_addr),
    .W0_clk(mem_0_16_W0_clk),
    .W0_data(mem_0_16_W0_data),
    .W0_en(mem_0_16_W0_en),
    .W0_mask(mem_0_16_W0_mask),
    .R0_addr(mem_0_16_R0_addr),
    .R0_clk(mem_0_16_R0_clk),
    .R0_data(mem_0_16_R0_data),
    .R0_en(mem_0_16_R0_en)
  );
  split_mem_0_ext mem_0_17 ( // @[:anonymous source@610.4]
    .W0_addr(mem_0_17_W0_addr),
    .W0_clk(mem_0_17_W0_clk),
    .W0_data(mem_0_17_W0_data),
    .W0_en(mem_0_17_W0_en),
    .W0_mask(mem_0_17_W0_mask),
    .R0_addr(mem_0_17_R0_addr),
    .R0_clk(mem_0_17_R0_clk),
    .R0_data(mem_0_17_R0_data),
    .R0_en(mem_0_17_R0_en)
  );
  split_mem_0_ext mem_0_18 ( // @[:anonymous source@611.4]
    .W0_addr(mem_0_18_W0_addr),
    .W0_clk(mem_0_18_W0_clk),
    .W0_data(mem_0_18_W0_data),
    .W0_en(mem_0_18_W0_en),
    .W0_mask(mem_0_18_W0_mask),
    .R0_addr(mem_0_18_R0_addr),
    .R0_clk(mem_0_18_R0_clk),
    .R0_data(mem_0_18_R0_data),
    .R0_en(mem_0_18_R0_en)
  );
  split_mem_0_ext mem_0_19 ( // @[:anonymous source@612.4]
    .W0_addr(mem_0_19_W0_addr),
    .W0_clk(mem_0_19_W0_clk),
    .W0_data(mem_0_19_W0_data),
    .W0_en(mem_0_19_W0_en),
    .W0_mask(mem_0_19_W0_mask),
    .R0_addr(mem_0_19_R0_addr),
    .R0_clk(mem_0_19_R0_clk),
    .R0_data(mem_0_19_R0_data),
    .R0_en(mem_0_19_R0_en)
  );
  split_mem_0_ext mem_0_20 ( // @[:anonymous source@613.4]
    .W0_addr(mem_0_20_W0_addr),
    .W0_clk(mem_0_20_W0_clk),
    .W0_data(mem_0_20_W0_data),
    .W0_en(mem_0_20_W0_en),
    .W0_mask(mem_0_20_W0_mask),
    .R0_addr(mem_0_20_R0_addr),
    .R0_clk(mem_0_20_R0_clk),
    .R0_data(mem_0_20_R0_data),
    .R0_en(mem_0_20_R0_en)
  );
  split_mem_0_ext mem_0_21 ( // @[:anonymous source@614.4]
    .W0_addr(mem_0_21_W0_addr),
    .W0_clk(mem_0_21_W0_clk),
    .W0_data(mem_0_21_W0_data),
    .W0_en(mem_0_21_W0_en),
    .W0_mask(mem_0_21_W0_mask),
    .R0_addr(mem_0_21_R0_addr),
    .R0_clk(mem_0_21_R0_clk),
    .R0_data(mem_0_21_R0_data),
    .R0_en(mem_0_21_R0_en)
  );
  split_mem_0_ext mem_0_22 ( // @[:anonymous source@615.4]
    .W0_addr(mem_0_22_W0_addr),
    .W0_clk(mem_0_22_W0_clk),
    .W0_data(mem_0_22_W0_data),
    .W0_en(mem_0_22_W0_en),
    .W0_mask(mem_0_22_W0_mask),
    .R0_addr(mem_0_22_R0_addr),
    .R0_clk(mem_0_22_R0_clk),
    .R0_data(mem_0_22_R0_data),
    .R0_en(mem_0_22_R0_en)
  );
  split_mem_0_ext mem_0_23 ( // @[:anonymous source@616.4]
    .W0_addr(mem_0_23_W0_addr),
    .W0_clk(mem_0_23_W0_clk),
    .W0_data(mem_0_23_W0_data),
    .W0_en(mem_0_23_W0_en),
    .W0_mask(mem_0_23_W0_mask),
    .R0_addr(mem_0_23_R0_addr),
    .R0_clk(mem_0_23_R0_clk),
    .R0_data(mem_0_23_R0_data),
    .R0_en(mem_0_23_R0_en)
  );
  split_mem_0_ext mem_0_24 ( // @[:anonymous source@617.4]
    .W0_addr(mem_0_24_W0_addr),
    .W0_clk(mem_0_24_W0_clk),
    .W0_data(mem_0_24_W0_data),
    .W0_en(mem_0_24_W0_en),
    .W0_mask(mem_0_24_W0_mask),
    .R0_addr(mem_0_24_R0_addr),
    .R0_clk(mem_0_24_R0_clk),
    .R0_data(mem_0_24_R0_data),
    .R0_en(mem_0_24_R0_en)
  );
  split_mem_0_ext mem_0_25 ( // @[:anonymous source@618.4]
    .W0_addr(mem_0_25_W0_addr),
    .W0_clk(mem_0_25_W0_clk),
    .W0_data(mem_0_25_W0_data),
    .W0_en(mem_0_25_W0_en),
    .W0_mask(mem_0_25_W0_mask),
    .R0_addr(mem_0_25_R0_addr),
    .R0_clk(mem_0_25_R0_clk),
    .R0_data(mem_0_25_R0_data),
    .R0_en(mem_0_25_R0_en)
  );
  split_mem_0_ext mem_0_26 ( // @[:anonymous source@619.4]
    .W0_addr(mem_0_26_W0_addr),
    .W0_clk(mem_0_26_W0_clk),
    .W0_data(mem_0_26_W0_data),
    .W0_en(mem_0_26_W0_en),
    .W0_mask(mem_0_26_W0_mask),
    .R0_addr(mem_0_26_R0_addr),
    .R0_clk(mem_0_26_R0_clk),
    .R0_data(mem_0_26_R0_data),
    .R0_en(mem_0_26_R0_en)
  );
  split_mem_0_ext mem_0_27 ( // @[:anonymous source@620.4]
    .W0_addr(mem_0_27_W0_addr),
    .W0_clk(mem_0_27_W0_clk),
    .W0_data(mem_0_27_W0_data),
    .W0_en(mem_0_27_W0_en),
    .W0_mask(mem_0_27_W0_mask),
    .R0_addr(mem_0_27_R0_addr),
    .R0_clk(mem_0_27_R0_clk),
    .R0_data(mem_0_27_R0_data),
    .R0_en(mem_0_27_R0_en)
  );
  split_mem_0_ext mem_0_28 ( // @[:anonymous source@621.4]
    .W0_addr(mem_0_28_W0_addr),
    .W0_clk(mem_0_28_W0_clk),
    .W0_data(mem_0_28_W0_data),
    .W0_en(mem_0_28_W0_en),
    .W0_mask(mem_0_28_W0_mask),
    .R0_addr(mem_0_28_R0_addr),
    .R0_clk(mem_0_28_R0_clk),
    .R0_data(mem_0_28_R0_data),
    .R0_en(mem_0_28_R0_en)
  );
  split_mem_0_ext mem_0_29 ( // @[:anonymous source@622.4]
    .W0_addr(mem_0_29_W0_addr),
    .W0_clk(mem_0_29_W0_clk),
    .W0_data(mem_0_29_W0_data),
    .W0_en(mem_0_29_W0_en),
    .W0_mask(mem_0_29_W0_mask),
    .R0_addr(mem_0_29_R0_addr),
    .R0_clk(mem_0_29_R0_clk),
    .R0_data(mem_0_29_R0_data),
    .R0_en(mem_0_29_R0_en)
  );
  split_mem_0_ext mem_0_30 ( // @[:anonymous source@623.4]
    .W0_addr(mem_0_30_W0_addr),
    .W0_clk(mem_0_30_W0_clk),
    .W0_data(mem_0_30_W0_data),
    .W0_en(mem_0_30_W0_en),
    .W0_mask(mem_0_30_W0_mask),
    .R0_addr(mem_0_30_R0_addr),
    .R0_clk(mem_0_30_R0_clk),
    .R0_data(mem_0_30_R0_data),
    .R0_en(mem_0_30_R0_en)
  );
  split_mem_0_ext mem_0_31 ( // @[:anonymous source@624.4]
    .W0_addr(mem_0_31_W0_addr),
    .W0_clk(mem_0_31_W0_clk),
    .W0_data(mem_0_31_W0_data),
    .W0_en(mem_0_31_W0_en),
    .W0_mask(mem_0_31_W0_mask),
    .R0_addr(mem_0_31_R0_addr),
    .R0_clk(mem_0_31_R0_clk),
    .R0_data(mem_0_31_R0_data),
    .R0_en(mem_0_31_R0_en)
  );
  split_mem_0_ext mem_0_32 ( // @[:anonymous source@625.4]
    .W0_addr(mem_0_32_W0_addr),
    .W0_clk(mem_0_32_W0_clk),
    .W0_data(mem_0_32_W0_data),
    .W0_en(mem_0_32_W0_en),
    .W0_mask(mem_0_32_W0_mask),
    .R0_addr(mem_0_32_R0_addr),
    .R0_clk(mem_0_32_R0_clk),
    .R0_data(mem_0_32_R0_data),
    .R0_en(mem_0_32_R0_en)
  );
  split_mem_0_ext mem_0_33 ( // @[:anonymous source@626.4]
    .W0_addr(mem_0_33_W0_addr),
    .W0_clk(mem_0_33_W0_clk),
    .W0_data(mem_0_33_W0_data),
    .W0_en(mem_0_33_W0_en),
    .W0_mask(mem_0_33_W0_mask),
    .R0_addr(mem_0_33_R0_addr),
    .R0_clk(mem_0_33_R0_clk),
    .R0_data(mem_0_33_R0_data),
    .R0_en(mem_0_33_R0_en)
  );
  split_mem_0_ext mem_0_34 ( // @[:anonymous source@627.4]
    .W0_addr(mem_0_34_W0_addr),
    .W0_clk(mem_0_34_W0_clk),
    .W0_data(mem_0_34_W0_data),
    .W0_en(mem_0_34_W0_en),
    .W0_mask(mem_0_34_W0_mask),
    .R0_addr(mem_0_34_R0_addr),
    .R0_clk(mem_0_34_R0_clk),
    .R0_data(mem_0_34_R0_data),
    .R0_en(mem_0_34_R0_en)
  );
  split_mem_0_ext mem_0_35 ( // @[:anonymous source@628.4]
    .W0_addr(mem_0_35_W0_addr),
    .W0_clk(mem_0_35_W0_clk),
    .W0_data(mem_0_35_W0_data),
    .W0_en(mem_0_35_W0_en),
    .W0_mask(mem_0_35_W0_mask),
    .R0_addr(mem_0_35_R0_addr),
    .R0_clk(mem_0_35_R0_clk),
    .R0_data(mem_0_35_R0_data),
    .R0_en(mem_0_35_R0_en)
  );
  split_mem_0_ext mem_0_36 ( // @[:anonymous source@629.4]
    .W0_addr(mem_0_36_W0_addr),
    .W0_clk(mem_0_36_W0_clk),
    .W0_data(mem_0_36_W0_data),
    .W0_en(mem_0_36_W0_en),
    .W0_mask(mem_0_36_W0_mask),
    .R0_addr(mem_0_36_R0_addr),
    .R0_clk(mem_0_36_R0_clk),
    .R0_data(mem_0_36_R0_data),
    .R0_en(mem_0_36_R0_en)
  );
  split_mem_0_ext mem_0_37 ( // @[:anonymous source@630.4]
    .W0_addr(mem_0_37_W0_addr),
    .W0_clk(mem_0_37_W0_clk),
    .W0_data(mem_0_37_W0_data),
    .W0_en(mem_0_37_W0_en),
    .W0_mask(mem_0_37_W0_mask),
    .R0_addr(mem_0_37_R0_addr),
    .R0_clk(mem_0_37_R0_clk),
    .R0_data(mem_0_37_R0_data),
    .R0_en(mem_0_37_R0_en)
  );
  split_mem_0_ext mem_0_38 ( // @[:anonymous source@631.4]
    .W0_addr(mem_0_38_W0_addr),
    .W0_clk(mem_0_38_W0_clk),
    .W0_data(mem_0_38_W0_data),
    .W0_en(mem_0_38_W0_en),
    .W0_mask(mem_0_38_W0_mask),
    .R0_addr(mem_0_38_R0_addr),
    .R0_clk(mem_0_38_R0_clk),
    .R0_data(mem_0_38_R0_data),
    .R0_en(mem_0_38_R0_en)
  );
  split_mem_0_ext mem_0_39 ( // @[:anonymous source@632.4]
    .W0_addr(mem_0_39_W0_addr),
    .W0_clk(mem_0_39_W0_clk),
    .W0_data(mem_0_39_W0_data),
    .W0_en(mem_0_39_W0_en),
    .W0_mask(mem_0_39_W0_mask),
    .R0_addr(mem_0_39_R0_addr),
    .R0_clk(mem_0_39_R0_clk),
    .R0_data(mem_0_39_R0_data),
    .R0_en(mem_0_39_R0_en)
  );
  split_mem_0_ext mem_0_40 ( // @[:anonymous source@633.4]
    .W0_addr(mem_0_40_W0_addr),
    .W0_clk(mem_0_40_W0_clk),
    .W0_data(mem_0_40_W0_data),
    .W0_en(mem_0_40_W0_en),
    .W0_mask(mem_0_40_W0_mask),
    .R0_addr(mem_0_40_R0_addr),
    .R0_clk(mem_0_40_R0_clk),
    .R0_data(mem_0_40_R0_data),
    .R0_en(mem_0_40_R0_en)
  );
  split_mem_0_ext mem_0_41 ( // @[:anonymous source@634.4]
    .W0_addr(mem_0_41_W0_addr),
    .W0_clk(mem_0_41_W0_clk),
    .W0_data(mem_0_41_W0_data),
    .W0_en(mem_0_41_W0_en),
    .W0_mask(mem_0_41_W0_mask),
    .R0_addr(mem_0_41_R0_addr),
    .R0_clk(mem_0_41_R0_clk),
    .R0_data(mem_0_41_R0_data),
    .R0_en(mem_0_41_R0_en)
  );
  split_mem_0_ext mem_0_42 ( // @[:anonymous source@635.4]
    .W0_addr(mem_0_42_W0_addr),
    .W0_clk(mem_0_42_W0_clk),
    .W0_data(mem_0_42_W0_data),
    .W0_en(mem_0_42_W0_en),
    .W0_mask(mem_0_42_W0_mask),
    .R0_addr(mem_0_42_R0_addr),
    .R0_clk(mem_0_42_R0_clk),
    .R0_data(mem_0_42_R0_data),
    .R0_en(mem_0_42_R0_en)
  );
  split_mem_0_ext mem_0_43 ( // @[:anonymous source@636.4]
    .W0_addr(mem_0_43_W0_addr),
    .W0_clk(mem_0_43_W0_clk),
    .W0_data(mem_0_43_W0_data),
    .W0_en(mem_0_43_W0_en),
    .W0_mask(mem_0_43_W0_mask),
    .R0_addr(mem_0_43_R0_addr),
    .R0_clk(mem_0_43_R0_clk),
    .R0_data(mem_0_43_R0_data),
    .R0_en(mem_0_43_R0_en)
  );
  split_mem_0_ext mem_0_44 ( // @[:anonymous source@637.4]
    .W0_addr(mem_0_44_W0_addr),
    .W0_clk(mem_0_44_W0_clk),
    .W0_data(mem_0_44_W0_data),
    .W0_en(mem_0_44_W0_en),
    .W0_mask(mem_0_44_W0_mask),
    .R0_addr(mem_0_44_R0_addr),
    .R0_clk(mem_0_44_R0_clk),
    .R0_data(mem_0_44_R0_data),
    .R0_en(mem_0_44_R0_en)
  );
  split_mem_0_ext mem_0_45 ( // @[:anonymous source@638.4]
    .W0_addr(mem_0_45_W0_addr),
    .W0_clk(mem_0_45_W0_clk),
    .W0_data(mem_0_45_W0_data),
    .W0_en(mem_0_45_W0_en),
    .W0_mask(mem_0_45_W0_mask),
    .R0_addr(mem_0_45_R0_addr),
    .R0_clk(mem_0_45_R0_clk),
    .R0_data(mem_0_45_R0_data),
    .R0_en(mem_0_45_R0_en)
  );
  split_mem_0_ext mem_0_46 ( // @[:anonymous source@639.4]
    .W0_addr(mem_0_46_W0_addr),
    .W0_clk(mem_0_46_W0_clk),
    .W0_data(mem_0_46_W0_data),
    .W0_en(mem_0_46_W0_en),
    .W0_mask(mem_0_46_W0_mask),
    .R0_addr(mem_0_46_R0_addr),
    .R0_clk(mem_0_46_R0_clk),
    .R0_data(mem_0_46_R0_data),
    .R0_en(mem_0_46_R0_en)
  );
  split_mem_0_ext mem_0_47 ( // @[:anonymous source@640.4]
    .W0_addr(mem_0_47_W0_addr),
    .W0_clk(mem_0_47_W0_clk),
    .W0_data(mem_0_47_W0_data),
    .W0_en(mem_0_47_W0_en),
    .W0_mask(mem_0_47_W0_mask),
    .R0_addr(mem_0_47_R0_addr),
    .R0_clk(mem_0_47_R0_clk),
    .R0_data(mem_0_47_R0_data),
    .R0_en(mem_0_47_R0_en)
  );
  split_mem_0_ext mem_0_48 ( // @[:anonymous source@641.4]
    .W0_addr(mem_0_48_W0_addr),
    .W0_clk(mem_0_48_W0_clk),
    .W0_data(mem_0_48_W0_data),
    .W0_en(mem_0_48_W0_en),
    .W0_mask(mem_0_48_W0_mask),
    .R0_addr(mem_0_48_R0_addr),
    .R0_clk(mem_0_48_R0_clk),
    .R0_data(mem_0_48_R0_data),
    .R0_en(mem_0_48_R0_en)
  );
  split_mem_0_ext mem_0_49 ( // @[:anonymous source@642.4]
    .W0_addr(mem_0_49_W0_addr),
    .W0_clk(mem_0_49_W0_clk),
    .W0_data(mem_0_49_W0_data),
    .W0_en(mem_0_49_W0_en),
    .W0_mask(mem_0_49_W0_mask),
    .R0_addr(mem_0_49_R0_addr),
    .R0_clk(mem_0_49_R0_clk),
    .R0_data(mem_0_49_R0_data),
    .R0_en(mem_0_49_R0_en)
  );
  split_mem_0_ext mem_0_50 ( // @[:anonymous source@643.4]
    .W0_addr(mem_0_50_W0_addr),
    .W0_clk(mem_0_50_W0_clk),
    .W0_data(mem_0_50_W0_data),
    .W0_en(mem_0_50_W0_en),
    .W0_mask(mem_0_50_W0_mask),
    .R0_addr(mem_0_50_R0_addr),
    .R0_clk(mem_0_50_R0_clk),
    .R0_data(mem_0_50_R0_data),
    .R0_en(mem_0_50_R0_en)
  );
  split_mem_0_ext mem_0_51 ( // @[:anonymous source@644.4]
    .W0_addr(mem_0_51_W0_addr),
    .W0_clk(mem_0_51_W0_clk),
    .W0_data(mem_0_51_W0_data),
    .W0_en(mem_0_51_W0_en),
    .W0_mask(mem_0_51_W0_mask),
    .R0_addr(mem_0_51_R0_addr),
    .R0_clk(mem_0_51_R0_clk),
    .R0_data(mem_0_51_R0_data),
    .R0_en(mem_0_51_R0_en)
  );
  split_mem_0_ext mem_0_52 ( // @[:anonymous source@645.4]
    .W0_addr(mem_0_52_W0_addr),
    .W0_clk(mem_0_52_W0_clk),
    .W0_data(mem_0_52_W0_data),
    .W0_en(mem_0_52_W0_en),
    .W0_mask(mem_0_52_W0_mask),
    .R0_addr(mem_0_52_R0_addr),
    .R0_clk(mem_0_52_R0_clk),
    .R0_data(mem_0_52_R0_data),
    .R0_en(mem_0_52_R0_en)
  );
  split_mem_0_ext mem_0_53 ( // @[:anonymous source@646.4]
    .W0_addr(mem_0_53_W0_addr),
    .W0_clk(mem_0_53_W0_clk),
    .W0_data(mem_0_53_W0_data),
    .W0_en(mem_0_53_W0_en),
    .W0_mask(mem_0_53_W0_mask),
    .R0_addr(mem_0_53_R0_addr),
    .R0_clk(mem_0_53_R0_clk),
    .R0_data(mem_0_53_R0_data),
    .R0_en(mem_0_53_R0_en)
  );
  split_mem_0_ext mem_0_54 ( // @[:anonymous source@647.4]
    .W0_addr(mem_0_54_W0_addr),
    .W0_clk(mem_0_54_W0_clk),
    .W0_data(mem_0_54_W0_data),
    .W0_en(mem_0_54_W0_en),
    .W0_mask(mem_0_54_W0_mask),
    .R0_addr(mem_0_54_R0_addr),
    .R0_clk(mem_0_54_R0_clk),
    .R0_data(mem_0_54_R0_data),
    .R0_en(mem_0_54_R0_en)
  );
  split_mem_0_ext mem_0_55 ( // @[:anonymous source@648.4]
    .W0_addr(mem_0_55_W0_addr),
    .W0_clk(mem_0_55_W0_clk),
    .W0_data(mem_0_55_W0_data),
    .W0_en(mem_0_55_W0_en),
    .W0_mask(mem_0_55_W0_mask),
    .R0_addr(mem_0_55_R0_addr),
    .R0_clk(mem_0_55_R0_clk),
    .R0_data(mem_0_55_R0_data),
    .R0_en(mem_0_55_R0_en)
  );
  split_mem_0_ext mem_0_56 ( // @[:anonymous source@649.4]
    .W0_addr(mem_0_56_W0_addr),
    .W0_clk(mem_0_56_W0_clk),
    .W0_data(mem_0_56_W0_data),
    .W0_en(mem_0_56_W0_en),
    .W0_mask(mem_0_56_W0_mask),
    .R0_addr(mem_0_56_R0_addr),
    .R0_clk(mem_0_56_R0_clk),
    .R0_data(mem_0_56_R0_data),
    .R0_en(mem_0_56_R0_en)
  );
  split_mem_0_ext mem_0_57 ( // @[:anonymous source@650.4]
    .W0_addr(mem_0_57_W0_addr),
    .W0_clk(mem_0_57_W0_clk),
    .W0_data(mem_0_57_W0_data),
    .W0_en(mem_0_57_W0_en),
    .W0_mask(mem_0_57_W0_mask),
    .R0_addr(mem_0_57_R0_addr),
    .R0_clk(mem_0_57_R0_clk),
    .R0_data(mem_0_57_R0_data),
    .R0_en(mem_0_57_R0_en)
  );
  split_mem_0_ext mem_0_58 ( // @[:anonymous source@651.4]
    .W0_addr(mem_0_58_W0_addr),
    .W0_clk(mem_0_58_W0_clk),
    .W0_data(mem_0_58_W0_data),
    .W0_en(mem_0_58_W0_en),
    .W0_mask(mem_0_58_W0_mask),
    .R0_addr(mem_0_58_R0_addr),
    .R0_clk(mem_0_58_R0_clk),
    .R0_data(mem_0_58_R0_data),
    .R0_en(mem_0_58_R0_en)
  );
  split_mem_0_ext mem_0_59 ( // @[:anonymous source@652.4]
    .W0_addr(mem_0_59_W0_addr),
    .W0_clk(mem_0_59_W0_clk),
    .W0_data(mem_0_59_W0_data),
    .W0_en(mem_0_59_W0_en),
    .W0_mask(mem_0_59_W0_mask),
    .R0_addr(mem_0_59_R0_addr),
    .R0_clk(mem_0_59_R0_clk),
    .R0_data(mem_0_59_R0_data),
    .R0_en(mem_0_59_R0_en)
  );
  split_mem_0_ext mem_0_60 ( // @[:anonymous source@653.4]
    .W0_addr(mem_0_60_W0_addr),
    .W0_clk(mem_0_60_W0_clk),
    .W0_data(mem_0_60_W0_data),
    .W0_en(mem_0_60_W0_en),
    .W0_mask(mem_0_60_W0_mask),
    .R0_addr(mem_0_60_R0_addr),
    .R0_clk(mem_0_60_R0_clk),
    .R0_data(mem_0_60_R0_data),
    .R0_en(mem_0_60_R0_en)
  );
  split_mem_0_ext mem_0_61 ( // @[:anonymous source@654.4]
    .W0_addr(mem_0_61_W0_addr),
    .W0_clk(mem_0_61_W0_clk),
    .W0_data(mem_0_61_W0_data),
    .W0_en(mem_0_61_W0_en),
    .W0_mask(mem_0_61_W0_mask),
    .R0_addr(mem_0_61_R0_addr),
    .R0_clk(mem_0_61_R0_clk),
    .R0_data(mem_0_61_R0_data),
    .R0_en(mem_0_61_R0_en)
  );
  split_mem_0_ext mem_0_62 ( // @[:anonymous source@655.4]
    .W0_addr(mem_0_62_W0_addr),
    .W0_clk(mem_0_62_W0_clk),
    .W0_data(mem_0_62_W0_data),
    .W0_en(mem_0_62_W0_en),
    .W0_mask(mem_0_62_W0_mask),
    .R0_addr(mem_0_62_R0_addr),
    .R0_clk(mem_0_62_R0_clk),
    .R0_data(mem_0_62_R0_data),
    .R0_en(mem_0_62_R0_en)
  );
  split_mem_0_ext mem_0_63 ( // @[:anonymous source@656.4]
    .W0_addr(mem_0_63_W0_addr),
    .W0_clk(mem_0_63_W0_clk),
    .W0_data(mem_0_63_W0_data),
    .W0_en(mem_0_63_W0_en),
    .W0_mask(mem_0_63_W0_mask),
    .R0_addr(mem_0_63_R0_addr),
    .R0_clk(mem_0_63_R0_clk),
    .R0_data(mem_0_63_R0_data),
    .R0_en(mem_0_63_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@979.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@983.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@987.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@991.4]
  assign R0_data_0_4 = mem_0_4_R0_data; // @[:anonymous source@995.4]
  assign R0_data_0_5 = mem_0_5_R0_data; // @[:anonymous source@999.4]
  assign R0_data_0_6 = mem_0_6_R0_data; // @[:anonymous source@1003.4]
  assign R0_data_0_7 = mem_0_7_R0_data; // @[:anonymous source@1007.4]
  assign R0_data_0_8 = mem_0_8_R0_data; // @[:anonymous source@1011.4]
  assign R0_data_0_9 = mem_0_9_R0_data; // @[:anonymous source@1015.4]
  assign R0_data_0_10 = mem_0_10_R0_data; // @[:anonymous source@1019.4]
  assign R0_data_0_11 = mem_0_11_R0_data; // @[:anonymous source@1023.4]
  assign R0_data_0_12 = mem_0_12_R0_data; // @[:anonymous source@1027.4]
  assign R0_data_0_13 = mem_0_13_R0_data; // @[:anonymous source@1031.4]
  assign R0_data_0_14 = mem_0_14_R0_data; // @[:anonymous source@1035.4]
  assign R0_data_0_15 = mem_0_15_R0_data; // @[:anonymous source@1039.4]
  assign R0_data_0_16 = mem_0_16_R0_data; // @[:anonymous source@1043.4]
  assign R0_data_0_17 = mem_0_17_R0_data; // @[:anonymous source@1047.4]
  assign R0_data_0_18 = mem_0_18_R0_data; // @[:anonymous source@1051.4]
  assign R0_data_0_19 = mem_0_19_R0_data; // @[:anonymous source@1055.4]
  assign R0_data_0_20 = mem_0_20_R0_data; // @[:anonymous source@1059.4]
  assign R0_data_0_21 = mem_0_21_R0_data; // @[:anonymous source@1063.4]
  assign R0_data_0_22 = mem_0_22_R0_data; // @[:anonymous source@1067.4]
  assign R0_data_0_23 = mem_0_23_R0_data; // @[:anonymous source@1071.4]
  assign R0_data_0_24 = mem_0_24_R0_data; // @[:anonymous source@1075.4]
  assign R0_data_0_25 = mem_0_25_R0_data; // @[:anonymous source@1079.4]
  assign R0_data_0_26 = mem_0_26_R0_data; // @[:anonymous source@1083.4]
  assign R0_data_0_27 = mem_0_27_R0_data; // @[:anonymous source@1087.4]
  assign R0_data_0_28 = mem_0_28_R0_data; // @[:anonymous source@1091.4]
  assign R0_data_0_29 = mem_0_29_R0_data; // @[:anonymous source@1095.4]
  assign R0_data_0_30 = mem_0_30_R0_data; // @[:anonymous source@1099.4]
  assign R0_data_0_31 = mem_0_31_R0_data; // @[:anonymous source@1103.4]
  assign R0_data_0_32 = mem_0_32_R0_data; // @[:anonymous source@1107.4]
  assign R0_data_0_33 = mem_0_33_R0_data; // @[:anonymous source@1111.4]
  assign R0_data_0_34 = mem_0_34_R0_data; // @[:anonymous source@1115.4]
  assign R0_data_0_35 = mem_0_35_R0_data; // @[:anonymous source@1119.4]
  assign R0_data_0_36 = mem_0_36_R0_data; // @[:anonymous source@1123.4]
  assign R0_data_0_37 = mem_0_37_R0_data; // @[:anonymous source@1127.4]
  assign R0_data_0_38 = mem_0_38_R0_data; // @[:anonymous source@1131.4]
  assign R0_data_0_39 = mem_0_39_R0_data; // @[:anonymous source@1135.4]
  assign R0_data_0_40 = mem_0_40_R0_data; // @[:anonymous source@1139.4]
  assign R0_data_0_41 = mem_0_41_R0_data; // @[:anonymous source@1143.4]
  assign R0_data_0_42 = mem_0_42_R0_data; // @[:anonymous source@1147.4]
  assign R0_data_0_43 = mem_0_43_R0_data; // @[:anonymous source@1151.4]
  assign R0_data_0_44 = mem_0_44_R0_data; // @[:anonymous source@1155.4]
  assign R0_data_0_45 = mem_0_45_R0_data; // @[:anonymous source@1159.4]
  assign R0_data_0_46 = mem_0_46_R0_data; // @[:anonymous source@1163.4]
  assign R0_data_0_47 = mem_0_47_R0_data; // @[:anonymous source@1167.4]
  assign R0_data_0_48 = mem_0_48_R0_data; // @[:anonymous source@1171.4]
  assign R0_data_0_49 = mem_0_49_R0_data; // @[:anonymous source@1175.4]
  assign R0_data_0_50 = mem_0_50_R0_data; // @[:anonymous source@1179.4]
  assign R0_data_0_51 = mem_0_51_R0_data; // @[:anonymous source@1183.4]
  assign R0_data_0_52 = mem_0_52_R0_data; // @[:anonymous source@1187.4]
  assign R0_data_0_53 = mem_0_53_R0_data; // @[:anonymous source@1191.4]
  assign R0_data_0_54 = mem_0_54_R0_data; // @[:anonymous source@1195.4]
  assign R0_data_0_55 = mem_0_55_R0_data; // @[:anonymous source@1199.4]
  assign R0_data_0_56 = mem_0_56_R0_data; // @[:anonymous source@1203.4]
  assign R0_data_0_57 = mem_0_57_R0_data; // @[:anonymous source@1207.4]
  assign R0_data_0_58 = mem_0_58_R0_data; // @[:anonymous source@1211.4]
  assign R0_data_0_59 = mem_0_59_R0_data; // @[:anonymous source@1215.4]
  assign R0_data_0_60 = mem_0_60_R0_data; // @[:anonymous source@1219.4]
  assign R0_data_0_61 = mem_0_61_R0_data; // @[:anonymous source@1223.4]
  assign R0_data_0_62 = mem_0_62_R0_data; // @[:anonymous source@1227.4]
  assign R0_data_0_63 = mem_0_63_R0_data; // @[:anonymous source@1231.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_2 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_3 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_4 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_5 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_6 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_7 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_8 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1233.4]
  assign _GEN_9 = {R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_10 = {R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_11 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_12 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_13 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_14 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_15 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_16 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_17 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1233.4]
  assign _GEN_18 = {R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_19 = {R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_20 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_21 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_22 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_23 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_24 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_25 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_26 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1233.4]
  assign _GEN_27 = {R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_28 = {R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_29 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_30 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_31 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_32 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_33 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_34 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_35 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1233.4]
  assign _GEN_36 = {R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_37 = {R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_38 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_39 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_40 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_41 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_42 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_43 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_44 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1233.4]
  assign _GEN_45 = {R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_46 = {R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_47 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_48 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_49 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_50 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_51 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_52 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_53 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1233.4]
  assign _GEN_54 = {R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_55 = {R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_56 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_57 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_58 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_59 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_60 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_61 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign R0_data_0 = {R0_data_0_63,R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1233.4]
  assign _GEN_62 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_63 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_64 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_65 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_66 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_67 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_68 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_69 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_70 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@1234.4]
  assign _GEN_71 = {R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_72 = {R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_73 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_74 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_75 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_76 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_77 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_78 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_79 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8}; // @[:anonymous source@1234.4]
  assign _GEN_80 = {R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_81 = {R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_82 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_83 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_84 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_85 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_86 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_87 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_88 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17}; // @[:anonymous source@1234.4]
  assign _GEN_89 = {R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_90 = {R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_91 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_92 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_93 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_94 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_95 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_96 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_97 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26}; // @[:anonymous source@1234.4]
  assign _GEN_98 = {R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_99 = {R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_100 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_101 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_102 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_103 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_104 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_105 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_106 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35}; // @[:anonymous source@1234.4]
  assign _GEN_107 = {R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_108 = {R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_109 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_110 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_111 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_112 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_113 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_114 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_115 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44}; // @[:anonymous source@1234.4]
  assign _GEN_116 = {R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_117 = {R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_118 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_119 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_120 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_121 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_122 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign _GEN_123 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53}; // @[:anonymous source@1234.4]
  assign R0_data = {R0_data_0_63,_GEN_61}; // @[:anonymous source@1234.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@658.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@657.4]
  assign mem_0_0_W0_data = W0_data[7:0]; // @[:anonymous source@659.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@661.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@660.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@978.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@977.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@980.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@663.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@662.4]
  assign mem_0_1_W0_data = W0_data[15:8]; // @[:anonymous source@664.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@666.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@665.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@982.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@981.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@984.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@668.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@667.4]
  assign mem_0_2_W0_data = W0_data[23:16]; // @[:anonymous source@669.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@671.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@670.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@986.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@985.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@988.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@673.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@672.4]
  assign mem_0_3_W0_data = W0_data[31:24]; // @[:anonymous source@674.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@676.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@675.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@990.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@989.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@992.4]
  assign mem_0_4_W0_addr = W0_addr; // @[:anonymous source@678.4]
  assign mem_0_4_W0_clk = W0_clk; // @[:anonymous source@677.4]
  assign mem_0_4_W0_data = W0_data[39:32]; // @[:anonymous source@679.4]
  assign mem_0_4_W0_en = W0_en; // @[:anonymous source@681.4]
  assign mem_0_4_W0_mask = W0_mask[4]; // @[:anonymous source@680.4]
  assign mem_0_4_R0_addr = R0_addr; // @[:anonymous source@994.4]
  assign mem_0_4_R0_clk = R0_clk; // @[:anonymous source@993.4]
  assign mem_0_4_R0_en = R0_en; // @[:anonymous source@996.4]
  assign mem_0_5_W0_addr = W0_addr; // @[:anonymous source@683.4]
  assign mem_0_5_W0_clk = W0_clk; // @[:anonymous source@682.4]
  assign mem_0_5_W0_data = W0_data[47:40]; // @[:anonymous source@684.4]
  assign mem_0_5_W0_en = W0_en; // @[:anonymous source@686.4]
  assign mem_0_5_W0_mask = W0_mask[5]; // @[:anonymous source@685.4]
  assign mem_0_5_R0_addr = R0_addr; // @[:anonymous source@998.4]
  assign mem_0_5_R0_clk = R0_clk; // @[:anonymous source@997.4]
  assign mem_0_5_R0_en = R0_en; // @[:anonymous source@1000.4]
  assign mem_0_6_W0_addr = W0_addr; // @[:anonymous source@688.4]
  assign mem_0_6_W0_clk = W0_clk; // @[:anonymous source@687.4]
  assign mem_0_6_W0_data = W0_data[55:48]; // @[:anonymous source@689.4]
  assign mem_0_6_W0_en = W0_en; // @[:anonymous source@691.4]
  assign mem_0_6_W0_mask = W0_mask[6]; // @[:anonymous source@690.4]
  assign mem_0_6_R0_addr = R0_addr; // @[:anonymous source@1002.4]
  assign mem_0_6_R0_clk = R0_clk; // @[:anonymous source@1001.4]
  assign mem_0_6_R0_en = R0_en; // @[:anonymous source@1004.4]
  assign mem_0_7_W0_addr = W0_addr; // @[:anonymous source@693.4]
  assign mem_0_7_W0_clk = W0_clk; // @[:anonymous source@692.4]
  assign mem_0_7_W0_data = W0_data[63:56]; // @[:anonymous source@694.4]
  assign mem_0_7_W0_en = W0_en; // @[:anonymous source@696.4]
  assign mem_0_7_W0_mask = W0_mask[7]; // @[:anonymous source@695.4]
  assign mem_0_7_R0_addr = R0_addr; // @[:anonymous source@1006.4]
  assign mem_0_7_R0_clk = R0_clk; // @[:anonymous source@1005.4]
  assign mem_0_7_R0_en = R0_en; // @[:anonymous source@1008.4]
  assign mem_0_8_W0_addr = W0_addr; // @[:anonymous source@698.4]
  assign mem_0_8_W0_clk = W0_clk; // @[:anonymous source@697.4]
  assign mem_0_8_W0_data = W0_data[71:64]; // @[:anonymous source@699.4]
  assign mem_0_8_W0_en = W0_en; // @[:anonymous source@701.4]
  assign mem_0_8_W0_mask = W0_mask[8]; // @[:anonymous source@700.4]
  assign mem_0_8_R0_addr = R0_addr; // @[:anonymous source@1010.4]
  assign mem_0_8_R0_clk = R0_clk; // @[:anonymous source@1009.4]
  assign mem_0_8_R0_en = R0_en; // @[:anonymous source@1012.4]
  assign mem_0_9_W0_addr = W0_addr; // @[:anonymous source@703.4]
  assign mem_0_9_W0_clk = W0_clk; // @[:anonymous source@702.4]
  assign mem_0_9_W0_data = W0_data[79:72]; // @[:anonymous source@704.4]
  assign mem_0_9_W0_en = W0_en; // @[:anonymous source@706.4]
  assign mem_0_9_W0_mask = W0_mask[9]; // @[:anonymous source@705.4]
  assign mem_0_9_R0_addr = R0_addr; // @[:anonymous source@1014.4]
  assign mem_0_9_R0_clk = R0_clk; // @[:anonymous source@1013.4]
  assign mem_0_9_R0_en = R0_en; // @[:anonymous source@1016.4]
  assign mem_0_10_W0_addr = W0_addr; // @[:anonymous source@708.4]
  assign mem_0_10_W0_clk = W0_clk; // @[:anonymous source@707.4]
  assign mem_0_10_W0_data = W0_data[87:80]; // @[:anonymous source@709.4]
  assign mem_0_10_W0_en = W0_en; // @[:anonymous source@711.4]
  assign mem_0_10_W0_mask = W0_mask[10]; // @[:anonymous source@710.4]
  assign mem_0_10_R0_addr = R0_addr; // @[:anonymous source@1018.4]
  assign mem_0_10_R0_clk = R0_clk; // @[:anonymous source@1017.4]
  assign mem_0_10_R0_en = R0_en; // @[:anonymous source@1020.4]
  assign mem_0_11_W0_addr = W0_addr; // @[:anonymous source@713.4]
  assign mem_0_11_W0_clk = W0_clk; // @[:anonymous source@712.4]
  assign mem_0_11_W0_data = W0_data[95:88]; // @[:anonymous source@714.4]
  assign mem_0_11_W0_en = W0_en; // @[:anonymous source@716.4]
  assign mem_0_11_W0_mask = W0_mask[11]; // @[:anonymous source@715.4]
  assign mem_0_11_R0_addr = R0_addr; // @[:anonymous source@1022.4]
  assign mem_0_11_R0_clk = R0_clk; // @[:anonymous source@1021.4]
  assign mem_0_11_R0_en = R0_en; // @[:anonymous source@1024.4]
  assign mem_0_12_W0_addr = W0_addr; // @[:anonymous source@718.4]
  assign mem_0_12_W0_clk = W0_clk; // @[:anonymous source@717.4]
  assign mem_0_12_W0_data = W0_data[103:96]; // @[:anonymous source@719.4]
  assign mem_0_12_W0_en = W0_en; // @[:anonymous source@721.4]
  assign mem_0_12_W0_mask = W0_mask[12]; // @[:anonymous source@720.4]
  assign mem_0_12_R0_addr = R0_addr; // @[:anonymous source@1026.4]
  assign mem_0_12_R0_clk = R0_clk; // @[:anonymous source@1025.4]
  assign mem_0_12_R0_en = R0_en; // @[:anonymous source@1028.4]
  assign mem_0_13_W0_addr = W0_addr; // @[:anonymous source@723.4]
  assign mem_0_13_W0_clk = W0_clk; // @[:anonymous source@722.4]
  assign mem_0_13_W0_data = W0_data[111:104]; // @[:anonymous source@724.4]
  assign mem_0_13_W0_en = W0_en; // @[:anonymous source@726.4]
  assign mem_0_13_W0_mask = W0_mask[13]; // @[:anonymous source@725.4]
  assign mem_0_13_R0_addr = R0_addr; // @[:anonymous source@1030.4]
  assign mem_0_13_R0_clk = R0_clk; // @[:anonymous source@1029.4]
  assign mem_0_13_R0_en = R0_en; // @[:anonymous source@1032.4]
  assign mem_0_14_W0_addr = W0_addr; // @[:anonymous source@728.4]
  assign mem_0_14_W0_clk = W0_clk; // @[:anonymous source@727.4]
  assign mem_0_14_W0_data = W0_data[119:112]; // @[:anonymous source@729.4]
  assign mem_0_14_W0_en = W0_en; // @[:anonymous source@731.4]
  assign mem_0_14_W0_mask = W0_mask[14]; // @[:anonymous source@730.4]
  assign mem_0_14_R0_addr = R0_addr; // @[:anonymous source@1034.4]
  assign mem_0_14_R0_clk = R0_clk; // @[:anonymous source@1033.4]
  assign mem_0_14_R0_en = R0_en; // @[:anonymous source@1036.4]
  assign mem_0_15_W0_addr = W0_addr; // @[:anonymous source@733.4]
  assign mem_0_15_W0_clk = W0_clk; // @[:anonymous source@732.4]
  assign mem_0_15_W0_data = W0_data[127:120]; // @[:anonymous source@734.4]
  assign mem_0_15_W0_en = W0_en; // @[:anonymous source@736.4]
  assign mem_0_15_W0_mask = W0_mask[15]; // @[:anonymous source@735.4]
  assign mem_0_15_R0_addr = R0_addr; // @[:anonymous source@1038.4]
  assign mem_0_15_R0_clk = R0_clk; // @[:anonymous source@1037.4]
  assign mem_0_15_R0_en = R0_en; // @[:anonymous source@1040.4]
  assign mem_0_16_W0_addr = W0_addr; // @[:anonymous source@738.4]
  assign mem_0_16_W0_clk = W0_clk; // @[:anonymous source@737.4]
  assign mem_0_16_W0_data = W0_data[135:128]; // @[:anonymous source@739.4]
  assign mem_0_16_W0_en = W0_en; // @[:anonymous source@741.4]
  assign mem_0_16_W0_mask = W0_mask[16]; // @[:anonymous source@740.4]
  assign mem_0_16_R0_addr = R0_addr; // @[:anonymous source@1042.4]
  assign mem_0_16_R0_clk = R0_clk; // @[:anonymous source@1041.4]
  assign mem_0_16_R0_en = R0_en; // @[:anonymous source@1044.4]
  assign mem_0_17_W0_addr = W0_addr; // @[:anonymous source@743.4]
  assign mem_0_17_W0_clk = W0_clk; // @[:anonymous source@742.4]
  assign mem_0_17_W0_data = W0_data[143:136]; // @[:anonymous source@744.4]
  assign mem_0_17_W0_en = W0_en; // @[:anonymous source@746.4]
  assign mem_0_17_W0_mask = W0_mask[17]; // @[:anonymous source@745.4]
  assign mem_0_17_R0_addr = R0_addr; // @[:anonymous source@1046.4]
  assign mem_0_17_R0_clk = R0_clk; // @[:anonymous source@1045.4]
  assign mem_0_17_R0_en = R0_en; // @[:anonymous source@1048.4]
  assign mem_0_18_W0_addr = W0_addr; // @[:anonymous source@748.4]
  assign mem_0_18_W0_clk = W0_clk; // @[:anonymous source@747.4]
  assign mem_0_18_W0_data = W0_data[151:144]; // @[:anonymous source@749.4]
  assign mem_0_18_W0_en = W0_en; // @[:anonymous source@751.4]
  assign mem_0_18_W0_mask = W0_mask[18]; // @[:anonymous source@750.4]
  assign mem_0_18_R0_addr = R0_addr; // @[:anonymous source@1050.4]
  assign mem_0_18_R0_clk = R0_clk; // @[:anonymous source@1049.4]
  assign mem_0_18_R0_en = R0_en; // @[:anonymous source@1052.4]
  assign mem_0_19_W0_addr = W0_addr; // @[:anonymous source@753.4]
  assign mem_0_19_W0_clk = W0_clk; // @[:anonymous source@752.4]
  assign mem_0_19_W0_data = W0_data[159:152]; // @[:anonymous source@754.4]
  assign mem_0_19_W0_en = W0_en; // @[:anonymous source@756.4]
  assign mem_0_19_W0_mask = W0_mask[19]; // @[:anonymous source@755.4]
  assign mem_0_19_R0_addr = R0_addr; // @[:anonymous source@1054.4]
  assign mem_0_19_R0_clk = R0_clk; // @[:anonymous source@1053.4]
  assign mem_0_19_R0_en = R0_en; // @[:anonymous source@1056.4]
  assign mem_0_20_W0_addr = W0_addr; // @[:anonymous source@758.4]
  assign mem_0_20_W0_clk = W0_clk; // @[:anonymous source@757.4]
  assign mem_0_20_W0_data = W0_data[167:160]; // @[:anonymous source@759.4]
  assign mem_0_20_W0_en = W0_en; // @[:anonymous source@761.4]
  assign mem_0_20_W0_mask = W0_mask[20]; // @[:anonymous source@760.4]
  assign mem_0_20_R0_addr = R0_addr; // @[:anonymous source@1058.4]
  assign mem_0_20_R0_clk = R0_clk; // @[:anonymous source@1057.4]
  assign mem_0_20_R0_en = R0_en; // @[:anonymous source@1060.4]
  assign mem_0_21_W0_addr = W0_addr; // @[:anonymous source@763.4]
  assign mem_0_21_W0_clk = W0_clk; // @[:anonymous source@762.4]
  assign mem_0_21_W0_data = W0_data[175:168]; // @[:anonymous source@764.4]
  assign mem_0_21_W0_en = W0_en; // @[:anonymous source@766.4]
  assign mem_0_21_W0_mask = W0_mask[21]; // @[:anonymous source@765.4]
  assign mem_0_21_R0_addr = R0_addr; // @[:anonymous source@1062.4]
  assign mem_0_21_R0_clk = R0_clk; // @[:anonymous source@1061.4]
  assign mem_0_21_R0_en = R0_en; // @[:anonymous source@1064.4]
  assign mem_0_22_W0_addr = W0_addr; // @[:anonymous source@768.4]
  assign mem_0_22_W0_clk = W0_clk; // @[:anonymous source@767.4]
  assign mem_0_22_W0_data = W0_data[183:176]; // @[:anonymous source@769.4]
  assign mem_0_22_W0_en = W0_en; // @[:anonymous source@771.4]
  assign mem_0_22_W0_mask = W0_mask[22]; // @[:anonymous source@770.4]
  assign mem_0_22_R0_addr = R0_addr; // @[:anonymous source@1066.4]
  assign mem_0_22_R0_clk = R0_clk; // @[:anonymous source@1065.4]
  assign mem_0_22_R0_en = R0_en; // @[:anonymous source@1068.4]
  assign mem_0_23_W0_addr = W0_addr; // @[:anonymous source@773.4]
  assign mem_0_23_W0_clk = W0_clk; // @[:anonymous source@772.4]
  assign mem_0_23_W0_data = W0_data[191:184]; // @[:anonymous source@774.4]
  assign mem_0_23_W0_en = W0_en; // @[:anonymous source@776.4]
  assign mem_0_23_W0_mask = W0_mask[23]; // @[:anonymous source@775.4]
  assign mem_0_23_R0_addr = R0_addr; // @[:anonymous source@1070.4]
  assign mem_0_23_R0_clk = R0_clk; // @[:anonymous source@1069.4]
  assign mem_0_23_R0_en = R0_en; // @[:anonymous source@1072.4]
  assign mem_0_24_W0_addr = W0_addr; // @[:anonymous source@778.4]
  assign mem_0_24_W0_clk = W0_clk; // @[:anonymous source@777.4]
  assign mem_0_24_W0_data = W0_data[199:192]; // @[:anonymous source@779.4]
  assign mem_0_24_W0_en = W0_en; // @[:anonymous source@781.4]
  assign mem_0_24_W0_mask = W0_mask[24]; // @[:anonymous source@780.4]
  assign mem_0_24_R0_addr = R0_addr; // @[:anonymous source@1074.4]
  assign mem_0_24_R0_clk = R0_clk; // @[:anonymous source@1073.4]
  assign mem_0_24_R0_en = R0_en; // @[:anonymous source@1076.4]
  assign mem_0_25_W0_addr = W0_addr; // @[:anonymous source@783.4]
  assign mem_0_25_W0_clk = W0_clk; // @[:anonymous source@782.4]
  assign mem_0_25_W0_data = W0_data[207:200]; // @[:anonymous source@784.4]
  assign mem_0_25_W0_en = W0_en; // @[:anonymous source@786.4]
  assign mem_0_25_W0_mask = W0_mask[25]; // @[:anonymous source@785.4]
  assign mem_0_25_R0_addr = R0_addr; // @[:anonymous source@1078.4]
  assign mem_0_25_R0_clk = R0_clk; // @[:anonymous source@1077.4]
  assign mem_0_25_R0_en = R0_en; // @[:anonymous source@1080.4]
  assign mem_0_26_W0_addr = W0_addr; // @[:anonymous source@788.4]
  assign mem_0_26_W0_clk = W0_clk; // @[:anonymous source@787.4]
  assign mem_0_26_W0_data = W0_data[215:208]; // @[:anonymous source@789.4]
  assign mem_0_26_W0_en = W0_en; // @[:anonymous source@791.4]
  assign mem_0_26_W0_mask = W0_mask[26]; // @[:anonymous source@790.4]
  assign mem_0_26_R0_addr = R0_addr; // @[:anonymous source@1082.4]
  assign mem_0_26_R0_clk = R0_clk; // @[:anonymous source@1081.4]
  assign mem_0_26_R0_en = R0_en; // @[:anonymous source@1084.4]
  assign mem_0_27_W0_addr = W0_addr; // @[:anonymous source@793.4]
  assign mem_0_27_W0_clk = W0_clk; // @[:anonymous source@792.4]
  assign mem_0_27_W0_data = W0_data[223:216]; // @[:anonymous source@794.4]
  assign mem_0_27_W0_en = W0_en; // @[:anonymous source@796.4]
  assign mem_0_27_W0_mask = W0_mask[27]; // @[:anonymous source@795.4]
  assign mem_0_27_R0_addr = R0_addr; // @[:anonymous source@1086.4]
  assign mem_0_27_R0_clk = R0_clk; // @[:anonymous source@1085.4]
  assign mem_0_27_R0_en = R0_en; // @[:anonymous source@1088.4]
  assign mem_0_28_W0_addr = W0_addr; // @[:anonymous source@798.4]
  assign mem_0_28_W0_clk = W0_clk; // @[:anonymous source@797.4]
  assign mem_0_28_W0_data = W0_data[231:224]; // @[:anonymous source@799.4]
  assign mem_0_28_W0_en = W0_en; // @[:anonymous source@801.4]
  assign mem_0_28_W0_mask = W0_mask[28]; // @[:anonymous source@800.4]
  assign mem_0_28_R0_addr = R0_addr; // @[:anonymous source@1090.4]
  assign mem_0_28_R0_clk = R0_clk; // @[:anonymous source@1089.4]
  assign mem_0_28_R0_en = R0_en; // @[:anonymous source@1092.4]
  assign mem_0_29_W0_addr = W0_addr; // @[:anonymous source@803.4]
  assign mem_0_29_W0_clk = W0_clk; // @[:anonymous source@802.4]
  assign mem_0_29_W0_data = W0_data[239:232]; // @[:anonymous source@804.4]
  assign mem_0_29_W0_en = W0_en; // @[:anonymous source@806.4]
  assign mem_0_29_W0_mask = W0_mask[29]; // @[:anonymous source@805.4]
  assign mem_0_29_R0_addr = R0_addr; // @[:anonymous source@1094.4]
  assign mem_0_29_R0_clk = R0_clk; // @[:anonymous source@1093.4]
  assign mem_0_29_R0_en = R0_en; // @[:anonymous source@1096.4]
  assign mem_0_30_W0_addr = W0_addr; // @[:anonymous source@808.4]
  assign mem_0_30_W0_clk = W0_clk; // @[:anonymous source@807.4]
  assign mem_0_30_W0_data = W0_data[247:240]; // @[:anonymous source@809.4]
  assign mem_0_30_W0_en = W0_en; // @[:anonymous source@811.4]
  assign mem_0_30_W0_mask = W0_mask[30]; // @[:anonymous source@810.4]
  assign mem_0_30_R0_addr = R0_addr; // @[:anonymous source@1098.4]
  assign mem_0_30_R0_clk = R0_clk; // @[:anonymous source@1097.4]
  assign mem_0_30_R0_en = R0_en; // @[:anonymous source@1100.4]
  assign mem_0_31_W0_addr = W0_addr; // @[:anonymous source@813.4]
  assign mem_0_31_W0_clk = W0_clk; // @[:anonymous source@812.4]
  assign mem_0_31_W0_data = W0_data[255:248]; // @[:anonymous source@814.4]
  assign mem_0_31_W0_en = W0_en; // @[:anonymous source@816.4]
  assign mem_0_31_W0_mask = W0_mask[31]; // @[:anonymous source@815.4]
  assign mem_0_31_R0_addr = R0_addr; // @[:anonymous source@1102.4]
  assign mem_0_31_R0_clk = R0_clk; // @[:anonymous source@1101.4]
  assign mem_0_31_R0_en = R0_en; // @[:anonymous source@1104.4]
  assign mem_0_32_W0_addr = W0_addr; // @[:anonymous source@818.4]
  assign mem_0_32_W0_clk = W0_clk; // @[:anonymous source@817.4]
  assign mem_0_32_W0_data = W0_data[263:256]; // @[:anonymous source@819.4]
  assign mem_0_32_W0_en = W0_en; // @[:anonymous source@821.4]
  assign mem_0_32_W0_mask = W0_mask[32]; // @[:anonymous source@820.4]
  assign mem_0_32_R0_addr = R0_addr; // @[:anonymous source@1106.4]
  assign mem_0_32_R0_clk = R0_clk; // @[:anonymous source@1105.4]
  assign mem_0_32_R0_en = R0_en; // @[:anonymous source@1108.4]
  assign mem_0_33_W0_addr = W0_addr; // @[:anonymous source@823.4]
  assign mem_0_33_W0_clk = W0_clk; // @[:anonymous source@822.4]
  assign mem_0_33_W0_data = W0_data[271:264]; // @[:anonymous source@824.4]
  assign mem_0_33_W0_en = W0_en; // @[:anonymous source@826.4]
  assign mem_0_33_W0_mask = W0_mask[33]; // @[:anonymous source@825.4]
  assign mem_0_33_R0_addr = R0_addr; // @[:anonymous source@1110.4]
  assign mem_0_33_R0_clk = R0_clk; // @[:anonymous source@1109.4]
  assign mem_0_33_R0_en = R0_en; // @[:anonymous source@1112.4]
  assign mem_0_34_W0_addr = W0_addr; // @[:anonymous source@828.4]
  assign mem_0_34_W0_clk = W0_clk; // @[:anonymous source@827.4]
  assign mem_0_34_W0_data = W0_data[279:272]; // @[:anonymous source@829.4]
  assign mem_0_34_W0_en = W0_en; // @[:anonymous source@831.4]
  assign mem_0_34_W0_mask = W0_mask[34]; // @[:anonymous source@830.4]
  assign mem_0_34_R0_addr = R0_addr; // @[:anonymous source@1114.4]
  assign mem_0_34_R0_clk = R0_clk; // @[:anonymous source@1113.4]
  assign mem_0_34_R0_en = R0_en; // @[:anonymous source@1116.4]
  assign mem_0_35_W0_addr = W0_addr; // @[:anonymous source@833.4]
  assign mem_0_35_W0_clk = W0_clk; // @[:anonymous source@832.4]
  assign mem_0_35_W0_data = W0_data[287:280]; // @[:anonymous source@834.4]
  assign mem_0_35_W0_en = W0_en; // @[:anonymous source@836.4]
  assign mem_0_35_W0_mask = W0_mask[35]; // @[:anonymous source@835.4]
  assign mem_0_35_R0_addr = R0_addr; // @[:anonymous source@1118.4]
  assign mem_0_35_R0_clk = R0_clk; // @[:anonymous source@1117.4]
  assign mem_0_35_R0_en = R0_en; // @[:anonymous source@1120.4]
  assign mem_0_36_W0_addr = W0_addr; // @[:anonymous source@838.4]
  assign mem_0_36_W0_clk = W0_clk; // @[:anonymous source@837.4]
  assign mem_0_36_W0_data = W0_data[295:288]; // @[:anonymous source@839.4]
  assign mem_0_36_W0_en = W0_en; // @[:anonymous source@841.4]
  assign mem_0_36_W0_mask = W0_mask[36]; // @[:anonymous source@840.4]
  assign mem_0_36_R0_addr = R0_addr; // @[:anonymous source@1122.4]
  assign mem_0_36_R0_clk = R0_clk; // @[:anonymous source@1121.4]
  assign mem_0_36_R0_en = R0_en; // @[:anonymous source@1124.4]
  assign mem_0_37_W0_addr = W0_addr; // @[:anonymous source@843.4]
  assign mem_0_37_W0_clk = W0_clk; // @[:anonymous source@842.4]
  assign mem_0_37_W0_data = W0_data[303:296]; // @[:anonymous source@844.4]
  assign mem_0_37_W0_en = W0_en; // @[:anonymous source@846.4]
  assign mem_0_37_W0_mask = W0_mask[37]; // @[:anonymous source@845.4]
  assign mem_0_37_R0_addr = R0_addr; // @[:anonymous source@1126.4]
  assign mem_0_37_R0_clk = R0_clk; // @[:anonymous source@1125.4]
  assign mem_0_37_R0_en = R0_en; // @[:anonymous source@1128.4]
  assign mem_0_38_W0_addr = W0_addr; // @[:anonymous source@848.4]
  assign mem_0_38_W0_clk = W0_clk; // @[:anonymous source@847.4]
  assign mem_0_38_W0_data = W0_data[311:304]; // @[:anonymous source@849.4]
  assign mem_0_38_W0_en = W0_en; // @[:anonymous source@851.4]
  assign mem_0_38_W0_mask = W0_mask[38]; // @[:anonymous source@850.4]
  assign mem_0_38_R0_addr = R0_addr; // @[:anonymous source@1130.4]
  assign mem_0_38_R0_clk = R0_clk; // @[:anonymous source@1129.4]
  assign mem_0_38_R0_en = R0_en; // @[:anonymous source@1132.4]
  assign mem_0_39_W0_addr = W0_addr; // @[:anonymous source@853.4]
  assign mem_0_39_W0_clk = W0_clk; // @[:anonymous source@852.4]
  assign mem_0_39_W0_data = W0_data[319:312]; // @[:anonymous source@854.4]
  assign mem_0_39_W0_en = W0_en; // @[:anonymous source@856.4]
  assign mem_0_39_W0_mask = W0_mask[39]; // @[:anonymous source@855.4]
  assign mem_0_39_R0_addr = R0_addr; // @[:anonymous source@1134.4]
  assign mem_0_39_R0_clk = R0_clk; // @[:anonymous source@1133.4]
  assign mem_0_39_R0_en = R0_en; // @[:anonymous source@1136.4]
  assign mem_0_40_W0_addr = W0_addr; // @[:anonymous source@858.4]
  assign mem_0_40_W0_clk = W0_clk; // @[:anonymous source@857.4]
  assign mem_0_40_W0_data = W0_data[327:320]; // @[:anonymous source@859.4]
  assign mem_0_40_W0_en = W0_en; // @[:anonymous source@861.4]
  assign mem_0_40_W0_mask = W0_mask[40]; // @[:anonymous source@860.4]
  assign mem_0_40_R0_addr = R0_addr; // @[:anonymous source@1138.4]
  assign mem_0_40_R0_clk = R0_clk; // @[:anonymous source@1137.4]
  assign mem_0_40_R0_en = R0_en; // @[:anonymous source@1140.4]
  assign mem_0_41_W0_addr = W0_addr; // @[:anonymous source@863.4]
  assign mem_0_41_W0_clk = W0_clk; // @[:anonymous source@862.4]
  assign mem_0_41_W0_data = W0_data[335:328]; // @[:anonymous source@864.4]
  assign mem_0_41_W0_en = W0_en; // @[:anonymous source@866.4]
  assign mem_0_41_W0_mask = W0_mask[41]; // @[:anonymous source@865.4]
  assign mem_0_41_R0_addr = R0_addr; // @[:anonymous source@1142.4]
  assign mem_0_41_R0_clk = R0_clk; // @[:anonymous source@1141.4]
  assign mem_0_41_R0_en = R0_en; // @[:anonymous source@1144.4]
  assign mem_0_42_W0_addr = W0_addr; // @[:anonymous source@868.4]
  assign mem_0_42_W0_clk = W0_clk; // @[:anonymous source@867.4]
  assign mem_0_42_W0_data = W0_data[343:336]; // @[:anonymous source@869.4]
  assign mem_0_42_W0_en = W0_en; // @[:anonymous source@871.4]
  assign mem_0_42_W0_mask = W0_mask[42]; // @[:anonymous source@870.4]
  assign mem_0_42_R0_addr = R0_addr; // @[:anonymous source@1146.4]
  assign mem_0_42_R0_clk = R0_clk; // @[:anonymous source@1145.4]
  assign mem_0_42_R0_en = R0_en; // @[:anonymous source@1148.4]
  assign mem_0_43_W0_addr = W0_addr; // @[:anonymous source@873.4]
  assign mem_0_43_W0_clk = W0_clk; // @[:anonymous source@872.4]
  assign mem_0_43_W0_data = W0_data[351:344]; // @[:anonymous source@874.4]
  assign mem_0_43_W0_en = W0_en; // @[:anonymous source@876.4]
  assign mem_0_43_W0_mask = W0_mask[43]; // @[:anonymous source@875.4]
  assign mem_0_43_R0_addr = R0_addr; // @[:anonymous source@1150.4]
  assign mem_0_43_R0_clk = R0_clk; // @[:anonymous source@1149.4]
  assign mem_0_43_R0_en = R0_en; // @[:anonymous source@1152.4]
  assign mem_0_44_W0_addr = W0_addr; // @[:anonymous source@878.4]
  assign mem_0_44_W0_clk = W0_clk; // @[:anonymous source@877.4]
  assign mem_0_44_W0_data = W0_data[359:352]; // @[:anonymous source@879.4]
  assign mem_0_44_W0_en = W0_en; // @[:anonymous source@881.4]
  assign mem_0_44_W0_mask = W0_mask[44]; // @[:anonymous source@880.4]
  assign mem_0_44_R0_addr = R0_addr; // @[:anonymous source@1154.4]
  assign mem_0_44_R0_clk = R0_clk; // @[:anonymous source@1153.4]
  assign mem_0_44_R0_en = R0_en; // @[:anonymous source@1156.4]
  assign mem_0_45_W0_addr = W0_addr; // @[:anonymous source@883.4]
  assign mem_0_45_W0_clk = W0_clk; // @[:anonymous source@882.4]
  assign mem_0_45_W0_data = W0_data[367:360]; // @[:anonymous source@884.4]
  assign mem_0_45_W0_en = W0_en; // @[:anonymous source@886.4]
  assign mem_0_45_W0_mask = W0_mask[45]; // @[:anonymous source@885.4]
  assign mem_0_45_R0_addr = R0_addr; // @[:anonymous source@1158.4]
  assign mem_0_45_R0_clk = R0_clk; // @[:anonymous source@1157.4]
  assign mem_0_45_R0_en = R0_en; // @[:anonymous source@1160.4]
  assign mem_0_46_W0_addr = W0_addr; // @[:anonymous source@888.4]
  assign mem_0_46_W0_clk = W0_clk; // @[:anonymous source@887.4]
  assign mem_0_46_W0_data = W0_data[375:368]; // @[:anonymous source@889.4]
  assign mem_0_46_W0_en = W0_en; // @[:anonymous source@891.4]
  assign mem_0_46_W0_mask = W0_mask[46]; // @[:anonymous source@890.4]
  assign mem_0_46_R0_addr = R0_addr; // @[:anonymous source@1162.4]
  assign mem_0_46_R0_clk = R0_clk; // @[:anonymous source@1161.4]
  assign mem_0_46_R0_en = R0_en; // @[:anonymous source@1164.4]
  assign mem_0_47_W0_addr = W0_addr; // @[:anonymous source@893.4]
  assign mem_0_47_W0_clk = W0_clk; // @[:anonymous source@892.4]
  assign mem_0_47_W0_data = W0_data[383:376]; // @[:anonymous source@894.4]
  assign mem_0_47_W0_en = W0_en; // @[:anonymous source@896.4]
  assign mem_0_47_W0_mask = W0_mask[47]; // @[:anonymous source@895.4]
  assign mem_0_47_R0_addr = R0_addr; // @[:anonymous source@1166.4]
  assign mem_0_47_R0_clk = R0_clk; // @[:anonymous source@1165.4]
  assign mem_0_47_R0_en = R0_en; // @[:anonymous source@1168.4]
  assign mem_0_48_W0_addr = W0_addr; // @[:anonymous source@898.4]
  assign mem_0_48_W0_clk = W0_clk; // @[:anonymous source@897.4]
  assign mem_0_48_W0_data = W0_data[391:384]; // @[:anonymous source@899.4]
  assign mem_0_48_W0_en = W0_en; // @[:anonymous source@901.4]
  assign mem_0_48_W0_mask = W0_mask[48]; // @[:anonymous source@900.4]
  assign mem_0_48_R0_addr = R0_addr; // @[:anonymous source@1170.4]
  assign mem_0_48_R0_clk = R0_clk; // @[:anonymous source@1169.4]
  assign mem_0_48_R0_en = R0_en; // @[:anonymous source@1172.4]
  assign mem_0_49_W0_addr = W0_addr; // @[:anonymous source@903.4]
  assign mem_0_49_W0_clk = W0_clk; // @[:anonymous source@902.4]
  assign mem_0_49_W0_data = W0_data[399:392]; // @[:anonymous source@904.4]
  assign mem_0_49_W0_en = W0_en; // @[:anonymous source@906.4]
  assign mem_0_49_W0_mask = W0_mask[49]; // @[:anonymous source@905.4]
  assign mem_0_49_R0_addr = R0_addr; // @[:anonymous source@1174.4]
  assign mem_0_49_R0_clk = R0_clk; // @[:anonymous source@1173.4]
  assign mem_0_49_R0_en = R0_en; // @[:anonymous source@1176.4]
  assign mem_0_50_W0_addr = W0_addr; // @[:anonymous source@908.4]
  assign mem_0_50_W0_clk = W0_clk; // @[:anonymous source@907.4]
  assign mem_0_50_W0_data = W0_data[407:400]; // @[:anonymous source@909.4]
  assign mem_0_50_W0_en = W0_en; // @[:anonymous source@911.4]
  assign mem_0_50_W0_mask = W0_mask[50]; // @[:anonymous source@910.4]
  assign mem_0_50_R0_addr = R0_addr; // @[:anonymous source@1178.4]
  assign mem_0_50_R0_clk = R0_clk; // @[:anonymous source@1177.4]
  assign mem_0_50_R0_en = R0_en; // @[:anonymous source@1180.4]
  assign mem_0_51_W0_addr = W0_addr; // @[:anonymous source@913.4]
  assign mem_0_51_W0_clk = W0_clk; // @[:anonymous source@912.4]
  assign mem_0_51_W0_data = W0_data[415:408]; // @[:anonymous source@914.4]
  assign mem_0_51_W0_en = W0_en; // @[:anonymous source@916.4]
  assign mem_0_51_W0_mask = W0_mask[51]; // @[:anonymous source@915.4]
  assign mem_0_51_R0_addr = R0_addr; // @[:anonymous source@1182.4]
  assign mem_0_51_R0_clk = R0_clk; // @[:anonymous source@1181.4]
  assign mem_0_51_R0_en = R0_en; // @[:anonymous source@1184.4]
  assign mem_0_52_W0_addr = W0_addr; // @[:anonymous source@918.4]
  assign mem_0_52_W0_clk = W0_clk; // @[:anonymous source@917.4]
  assign mem_0_52_W0_data = W0_data[423:416]; // @[:anonymous source@919.4]
  assign mem_0_52_W0_en = W0_en; // @[:anonymous source@921.4]
  assign mem_0_52_W0_mask = W0_mask[52]; // @[:anonymous source@920.4]
  assign mem_0_52_R0_addr = R0_addr; // @[:anonymous source@1186.4]
  assign mem_0_52_R0_clk = R0_clk; // @[:anonymous source@1185.4]
  assign mem_0_52_R0_en = R0_en; // @[:anonymous source@1188.4]
  assign mem_0_53_W0_addr = W0_addr; // @[:anonymous source@923.4]
  assign mem_0_53_W0_clk = W0_clk; // @[:anonymous source@922.4]
  assign mem_0_53_W0_data = W0_data[431:424]; // @[:anonymous source@924.4]
  assign mem_0_53_W0_en = W0_en; // @[:anonymous source@926.4]
  assign mem_0_53_W0_mask = W0_mask[53]; // @[:anonymous source@925.4]
  assign mem_0_53_R0_addr = R0_addr; // @[:anonymous source@1190.4]
  assign mem_0_53_R0_clk = R0_clk; // @[:anonymous source@1189.4]
  assign mem_0_53_R0_en = R0_en; // @[:anonymous source@1192.4]
  assign mem_0_54_W0_addr = W0_addr; // @[:anonymous source@928.4]
  assign mem_0_54_W0_clk = W0_clk; // @[:anonymous source@927.4]
  assign mem_0_54_W0_data = W0_data[439:432]; // @[:anonymous source@929.4]
  assign mem_0_54_W0_en = W0_en; // @[:anonymous source@931.4]
  assign mem_0_54_W0_mask = W0_mask[54]; // @[:anonymous source@930.4]
  assign mem_0_54_R0_addr = R0_addr; // @[:anonymous source@1194.4]
  assign mem_0_54_R0_clk = R0_clk; // @[:anonymous source@1193.4]
  assign mem_0_54_R0_en = R0_en; // @[:anonymous source@1196.4]
  assign mem_0_55_W0_addr = W0_addr; // @[:anonymous source@933.4]
  assign mem_0_55_W0_clk = W0_clk; // @[:anonymous source@932.4]
  assign mem_0_55_W0_data = W0_data[447:440]; // @[:anonymous source@934.4]
  assign mem_0_55_W0_en = W0_en; // @[:anonymous source@936.4]
  assign mem_0_55_W0_mask = W0_mask[55]; // @[:anonymous source@935.4]
  assign mem_0_55_R0_addr = R0_addr; // @[:anonymous source@1198.4]
  assign mem_0_55_R0_clk = R0_clk; // @[:anonymous source@1197.4]
  assign mem_0_55_R0_en = R0_en; // @[:anonymous source@1200.4]
  assign mem_0_56_W0_addr = W0_addr; // @[:anonymous source@938.4]
  assign mem_0_56_W0_clk = W0_clk; // @[:anonymous source@937.4]
  assign mem_0_56_W0_data = W0_data[455:448]; // @[:anonymous source@939.4]
  assign mem_0_56_W0_en = W0_en; // @[:anonymous source@941.4]
  assign mem_0_56_W0_mask = W0_mask[56]; // @[:anonymous source@940.4]
  assign mem_0_56_R0_addr = R0_addr; // @[:anonymous source@1202.4]
  assign mem_0_56_R0_clk = R0_clk; // @[:anonymous source@1201.4]
  assign mem_0_56_R0_en = R0_en; // @[:anonymous source@1204.4]
  assign mem_0_57_W0_addr = W0_addr; // @[:anonymous source@943.4]
  assign mem_0_57_W0_clk = W0_clk; // @[:anonymous source@942.4]
  assign mem_0_57_W0_data = W0_data[463:456]; // @[:anonymous source@944.4]
  assign mem_0_57_W0_en = W0_en; // @[:anonymous source@946.4]
  assign mem_0_57_W0_mask = W0_mask[57]; // @[:anonymous source@945.4]
  assign mem_0_57_R0_addr = R0_addr; // @[:anonymous source@1206.4]
  assign mem_0_57_R0_clk = R0_clk; // @[:anonymous source@1205.4]
  assign mem_0_57_R0_en = R0_en; // @[:anonymous source@1208.4]
  assign mem_0_58_W0_addr = W0_addr; // @[:anonymous source@948.4]
  assign mem_0_58_W0_clk = W0_clk; // @[:anonymous source@947.4]
  assign mem_0_58_W0_data = W0_data[471:464]; // @[:anonymous source@949.4]
  assign mem_0_58_W0_en = W0_en; // @[:anonymous source@951.4]
  assign mem_0_58_W0_mask = W0_mask[58]; // @[:anonymous source@950.4]
  assign mem_0_58_R0_addr = R0_addr; // @[:anonymous source@1210.4]
  assign mem_0_58_R0_clk = R0_clk; // @[:anonymous source@1209.4]
  assign mem_0_58_R0_en = R0_en; // @[:anonymous source@1212.4]
  assign mem_0_59_W0_addr = W0_addr; // @[:anonymous source@953.4]
  assign mem_0_59_W0_clk = W0_clk; // @[:anonymous source@952.4]
  assign mem_0_59_W0_data = W0_data[479:472]; // @[:anonymous source@954.4]
  assign mem_0_59_W0_en = W0_en; // @[:anonymous source@956.4]
  assign mem_0_59_W0_mask = W0_mask[59]; // @[:anonymous source@955.4]
  assign mem_0_59_R0_addr = R0_addr; // @[:anonymous source@1214.4]
  assign mem_0_59_R0_clk = R0_clk; // @[:anonymous source@1213.4]
  assign mem_0_59_R0_en = R0_en; // @[:anonymous source@1216.4]
  assign mem_0_60_W0_addr = W0_addr; // @[:anonymous source@958.4]
  assign mem_0_60_W0_clk = W0_clk; // @[:anonymous source@957.4]
  assign mem_0_60_W0_data = W0_data[487:480]; // @[:anonymous source@959.4]
  assign mem_0_60_W0_en = W0_en; // @[:anonymous source@961.4]
  assign mem_0_60_W0_mask = W0_mask[60]; // @[:anonymous source@960.4]
  assign mem_0_60_R0_addr = R0_addr; // @[:anonymous source@1218.4]
  assign mem_0_60_R0_clk = R0_clk; // @[:anonymous source@1217.4]
  assign mem_0_60_R0_en = R0_en; // @[:anonymous source@1220.4]
  assign mem_0_61_W0_addr = W0_addr; // @[:anonymous source@963.4]
  assign mem_0_61_W0_clk = W0_clk; // @[:anonymous source@962.4]
  assign mem_0_61_W0_data = W0_data[495:488]; // @[:anonymous source@964.4]
  assign mem_0_61_W0_en = W0_en; // @[:anonymous source@966.4]
  assign mem_0_61_W0_mask = W0_mask[61]; // @[:anonymous source@965.4]
  assign mem_0_61_R0_addr = R0_addr; // @[:anonymous source@1222.4]
  assign mem_0_61_R0_clk = R0_clk; // @[:anonymous source@1221.4]
  assign mem_0_61_R0_en = R0_en; // @[:anonymous source@1224.4]
  assign mem_0_62_W0_addr = W0_addr; // @[:anonymous source@968.4]
  assign mem_0_62_W0_clk = W0_clk; // @[:anonymous source@967.4]
  assign mem_0_62_W0_data = W0_data[503:496]; // @[:anonymous source@969.4]
  assign mem_0_62_W0_en = W0_en; // @[:anonymous source@971.4]
  assign mem_0_62_W0_mask = W0_mask[62]; // @[:anonymous source@970.4]
  assign mem_0_62_R0_addr = R0_addr; // @[:anonymous source@1226.4]
  assign mem_0_62_R0_clk = R0_clk; // @[:anonymous source@1225.4]
  assign mem_0_62_R0_en = R0_en; // @[:anonymous source@1228.4]
  assign mem_0_63_W0_addr = W0_addr; // @[:anonymous source@973.4]
  assign mem_0_63_W0_clk = W0_clk; // @[:anonymous source@972.4]
  assign mem_0_63_W0_data = W0_data[511:504]; // @[:anonymous source@974.4]
  assign mem_0_63_W0_en = W0_en; // @[:anonymous source@976.4]
  assign mem_0_63_W0_mask = W0_mask[63]; // @[:anonymous source@975.4]
  assign mem_0_63_R0_addr = R0_addr; // @[:anonymous source@1230.4]
  assign mem_0_63_R0_clk = R0_clk; // @[:anonymous source@1229.4]
  assign mem_0_63_R0_en = R0_en; // @[:anonymous source@1232.4]
endmodule
module tag_array_0_ext( // @[:anonymous source@1236.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@1237.4]
  input         RW0_clk, // @[:anonymous source@1238.4]
  input  [83:0] RW0_wdata, // @[:anonymous source@1239.4]
  output [83:0] RW0_rdata, // @[:anonymous source@1240.4]
  input         RW0_en, // @[:anonymous source@1241.4]
  input         RW0_wmode, // @[:anonymous source@1242.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@1243.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@1245.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@1245.4]
  wire [20:0] mem_0_0_RW0_wdata; // @[:anonymous source@1245.4]
  wire [20:0] mem_0_0_RW0_rdata; // @[:anonymous source@1245.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@1245.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@1245.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@1245.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@1246.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@1246.4]
  wire [20:0] mem_0_1_RW0_wdata; // @[:anonymous source@1246.4]
  wire [20:0] mem_0_1_RW0_rdata; // @[:anonymous source@1246.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@1246.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@1246.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@1246.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@1247.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@1247.4]
  wire [20:0] mem_0_2_RW0_wdata; // @[:anonymous source@1247.4]
  wire [20:0] mem_0_2_RW0_rdata; // @[:anonymous source@1247.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@1247.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@1247.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@1247.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@1248.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@1248.4]
  wire [20:0] mem_0_3_RW0_wdata; // @[:anonymous source@1248.4]
  wire [20:0] mem_0_3_RW0_rdata; // @[:anonymous source@1248.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@1248.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@1248.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@1248.4]
  wire [20:0] RW0_rdata_0_0; // @[:anonymous source@1251.4]
  wire [20:0] RW0_rdata_0_1; // @[:anonymous source@1258.4]
  wire [20:0] RW0_rdata_0_2; // @[:anonymous source@1265.4]
  wire [20:0] RW0_rdata_0_3; // @[:anonymous source@1272.4]
  wire [41:0] _GEN_0; // @[:anonymous source@1277.4]
  wire [62:0] _GEN_1; // @[:anonymous source@1277.4]
  wire [83:0] RW0_rdata_0; // @[:anonymous source@1277.4]
  wire [41:0] _GEN_2; // @[:anonymous source@1278.4]
  wire [62:0] _GEN_3; // @[:anonymous source@1278.4]
  split_tag_array_0_ext mem_0_0 ( // @[:anonymous source@1245.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 ( // @[:anonymous source@1246.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 ( // @[:anonymous source@1247.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 ( // @[:anonymous source@1248.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@1251.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@1258.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@1265.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@1272.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1277.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1277.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1277.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1278.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1278.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@1278.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@1250.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@1249.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[20:0]; // @[:anonymous source@1252.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@1255.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@1254.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@1253.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@1257.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@1256.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[41:21]; // @[:anonymous source@1259.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@1262.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@1261.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@1260.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@1264.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@1263.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[62:42]; // @[:anonymous source@1266.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@1269.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@1268.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@1267.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@1271.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@1270.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[83:63]; // @[:anonymous source@1273.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@1276.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@1275.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@1274.4]
endmodule
module data_arrays_0_0_ext( // @[:anonymous source@1280.2]
  input  [7:0]   RW0_addr, // @[:anonymous source@1281.4]
  input          RW0_clk, // @[:anonymous source@1282.4]
  input  [127:0] RW0_wdata, // @[:anonymous source@1283.4]
  output [127:0] RW0_rdata, // @[:anonymous source@1284.4]
  input          RW0_en, // @[:anonymous source@1285.4]
  input          RW0_wmode, // @[:anonymous source@1286.4]
  input  [3:0]   RW0_wmask // @[:anonymous source@1287.4]
);
  wire [7:0] mem_0_0_RW0_addr; // @[:anonymous source@1289.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@1289.4]
  wire [31:0] mem_0_0_RW0_wdata; // @[:anonymous source@1289.4]
  wire [31:0] mem_0_0_RW0_rdata; // @[:anonymous source@1289.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@1289.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@1289.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@1289.4]
  wire [7:0] mem_0_1_RW0_addr; // @[:anonymous source@1290.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@1290.4]
  wire [31:0] mem_0_1_RW0_wdata; // @[:anonymous source@1290.4]
  wire [31:0] mem_0_1_RW0_rdata; // @[:anonymous source@1290.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@1290.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@1290.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@1290.4]
  wire [7:0] mem_0_2_RW0_addr; // @[:anonymous source@1291.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@1291.4]
  wire [31:0] mem_0_2_RW0_wdata; // @[:anonymous source@1291.4]
  wire [31:0] mem_0_2_RW0_rdata; // @[:anonymous source@1291.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@1291.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@1291.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@1291.4]
  wire [7:0] mem_0_3_RW0_addr; // @[:anonymous source@1292.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@1292.4]
  wire [31:0] mem_0_3_RW0_wdata; // @[:anonymous source@1292.4]
  wire [31:0] mem_0_3_RW0_rdata; // @[:anonymous source@1292.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@1292.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@1292.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@1292.4]
  wire [31:0] RW0_rdata_0_0; // @[:anonymous source@1295.4]
  wire [31:0] RW0_rdata_0_1; // @[:anonymous source@1302.4]
  wire [31:0] RW0_rdata_0_2; // @[:anonymous source@1309.4]
  wire [31:0] RW0_rdata_0_3; // @[:anonymous source@1316.4]
  wire [63:0] _GEN_0; // @[:anonymous source@1321.4]
  wire [95:0] _GEN_1; // @[:anonymous source@1321.4]
  wire [127:0] RW0_rdata_0; // @[:anonymous source@1321.4]
  wire [63:0] _GEN_2; // @[:anonymous source@1322.4]
  wire [95:0] _GEN_3; // @[:anonymous source@1322.4]
  split_data_arrays_0_0_ext mem_0_0 ( // @[:anonymous source@1289.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_1 ( // @[:anonymous source@1290.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_2 ( // @[:anonymous source@1291.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_3 ( // @[:anonymous source@1292.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@1295.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@1302.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@1309.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@1316.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1321.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1321.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1321.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1322.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@1322.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@1322.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@1294.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@1293.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[31:0]; // @[:anonymous source@1296.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@1299.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@1298.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@1297.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@1301.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@1300.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[63:32]; // @[:anonymous source@1303.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@1306.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@1305.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@1304.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@1308.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@1307.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[95:64]; // @[:anonymous source@1310.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@1313.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@1312.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@1311.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@1315.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@1314.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[127:96]; // @[:anonymous source@1317.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@1320.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@1319.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@1318.4]
endmodule
module l2_tlb_ram_ext( // @[:anonymous source@1324.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1325.4]
  input         RW0_clk, // @[:anonymous source@1326.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@1327.4]
  output [43:0] RW0_rdata, // @[:anonymous source@1328.4]
  input         RW0_en, // @[:anonymous source@1329.4]
  input         RW0_wmode // @[:anonymous source@1330.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@1332.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@1332.4]
  wire [43:0] mem_0_0_RW0_wdata; // @[:anonymous source@1332.4]
  wire [43:0] mem_0_0_RW0_rdata; // @[:anonymous source@1332.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@1332.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@1332.4]
  wire [43:0] RW0_rdata_0_0; // @[:anonymous source@1335.4]
  wire [43:0] RW0_rdata_0; // @[:anonymous source@1339.4]
  split_l2_tlb_ram_ext mem_0_0 ( // @[:anonymous source@1332.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@1335.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@1339.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@1340.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@1334.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@1333.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@1336.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@1338.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@1337.4]
endmodule
module split_cc_dir_ext( // @[:anonymous source@1342.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1343.4]
  input         RW0_clk, // @[:anonymous source@1344.4]
  input  [15:0] RW0_wdata, // @[:anonymous source@1345.4]
  output [15:0] RW0_rdata, // @[:anonymous source@1346.4]
  input         RW0_en, // @[:anonymous source@1347.4]
  input         RW0_wmode, // @[:anonymous source@1348.4]
  input         RW0_wmask // @[:anonymous source@1349.4]
);
  reg [15:0] ram [0:1023]; // @[:anonymous source@1351.4]
  reg [31:0] _RAND_0;
  wire [15:0] ram_RW_0_r_data; // @[:anonymous source@1351.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@1351.4]
  wire [15:0] ram_RW_0_w_data; // @[:anonymous source@1351.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@1351.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1351.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1351.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1351.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1363.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1351.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_cc_banks_0_ext( // @[:anonymous source@1366.2]
  input  [12:0] RW0_addr, // @[:anonymous source@1367.4]
  input         RW0_clk, // @[:anonymous source@1368.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@1369.4]
  output [63:0] RW0_rdata, // @[:anonymous source@1370.4]
  input         RW0_en, // @[:anonymous source@1371.4]
  input         RW0_wmode // @[:anonymous source@1372.4]
);
  reg [63:0] ram [0:8191]; // @[:anonymous source@1374.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@1374.4]
  wire [12:0] ram_RW_0_r_addr; // @[:anonymous source@1374.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@1374.4]
  wire [12:0] ram_RW_0_w_addr; // @[:anonymous source@1374.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1374.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1374.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [12:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1374.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1386.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1374.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_data_arrays_0_ext( // @[:anonymous source@1389.2]
  input  [7:0] RW0_addr, // @[:anonymous source@1390.4]
  input        RW0_clk, // @[:anonymous source@1391.4]
  input  [7:0] RW0_wdata, // @[:anonymous source@1392.4]
  output [7:0] RW0_rdata, // @[:anonymous source@1393.4]
  input        RW0_en, // @[:anonymous source@1394.4]
  input        RW0_wmode, // @[:anonymous source@1395.4]
  input        RW0_wmask // @[:anonymous source@1396.4]
);
  reg [7:0] ram [0:255]; // @[:anonymous source@1398.4]
  reg [31:0] _RAND_0;
  wire [7:0] ram_RW_0_r_data; // @[:anonymous source@1398.4]
  wire [7:0] ram_RW_0_r_addr; // @[:anonymous source@1398.4]
  wire [7:0] ram_RW_0_w_data; // @[:anonymous source@1398.4]
  wire [7:0] ram_RW_0_w_addr; // @[:anonymous source@1398.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1398.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1398.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1398.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1410.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1398.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_tag_array_ext( // @[:anonymous source@1413.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@1414.4]
  input         RW0_clk, // @[:anonymous source@1415.4]
  input  [21:0] RW0_wdata, // @[:anonymous source@1416.4]
  output [21:0] RW0_rdata, // @[:anonymous source@1417.4]
  input         RW0_en, // @[:anonymous source@1418.4]
  input         RW0_wmode, // @[:anonymous source@1419.4]
  input         RW0_wmask // @[:anonymous source@1420.4]
);
  reg [21:0] ram [0:63]; // @[:anonymous source@1422.4]
  reg [31:0] _RAND_0;
  wire [21:0] ram_RW_0_r_data; // @[:anonymous source@1422.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@1422.4]
  wire [21:0] ram_RW_0_w_data; // @[:anonymous source@1422.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@1422.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1422.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1422.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1422.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1434.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1422.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_mem_ext( // @[:anonymous source@1437.2]
  input  [11:0] W0_addr, // @[:anonymous source@1438.4]
  input         W0_clk, // @[:anonymous source@1439.4]
  input  [7:0]  W0_data, // @[:anonymous source@1440.4]
  input         W0_en, // @[:anonymous source@1441.4]
  input         W0_mask, // @[:anonymous source@1442.4]
  input  [11:0] R0_addr, // @[:anonymous source@1443.4]
  input         R0_clk, // @[:anonymous source@1444.4]
  output [7:0]  R0_data, // @[:anonymous source@1445.4]
  input         R0_en // @[:anonymous source@1446.4]
);
  reg [7:0] ram [0:4095]; // @[:anonymous source@1448.4]
  reg [31:0] _RAND_0;
  wire [7:0] ram_R_0_data; // @[:anonymous source@1448.4]
  wire [11:0] ram_R_0_addr; // @[:anonymous source@1448.4]
  wire [7:0] ram_W_0_data; // @[:anonymous source@1448.4]
  wire [11:0] ram_W_0_addr; // @[:anonymous source@1448.4]
  wire  ram_W_0_mask; // @[:anonymous source@1448.4]
  wire  ram_W_0_en; // @[:anonymous source@1448.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [11:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1448.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1459.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[11:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1448.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_mem_0_ext( // @[:anonymous source@1466.2]
  input  [9:0] W0_addr, // @[:anonymous source@1467.4]
  input        W0_clk, // @[:anonymous source@1468.4]
  input  [7:0] W0_data, // @[:anonymous source@1469.4]
  input        W0_en, // @[:anonymous source@1470.4]
  input        W0_mask, // @[:anonymous source@1471.4]
  input  [9:0] R0_addr, // @[:anonymous source@1472.4]
  input        R0_clk, // @[:anonymous source@1473.4]
  output [7:0] R0_data, // @[:anonymous source@1474.4]
  input        R0_en // @[:anonymous source@1475.4]
);
  reg [7:0] ram [0:1023]; // @[:anonymous source@1477.4]
  reg [31:0] _RAND_0;
  wire [7:0] ram_R_0_data; // @[:anonymous source@1477.4]
  wire [9:0] ram_R_0_addr; // @[:anonymous source@1477.4]
  wire [7:0] ram_W_0_data; // @[:anonymous source@1477.4]
  wire [9:0] ram_W_0_addr; // @[:anonymous source@1477.4]
  wire  ram_W_0_mask; // @[:anonymous source@1477.4]
  wire  ram_W_0_en; // @[:anonymous source@1477.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1477.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1488.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1477.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_tag_array_0_ext( // @[:anonymous source@1495.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@1496.4]
  input         RW0_clk, // @[:anonymous source@1497.4]
  input  [20:0] RW0_wdata, // @[:anonymous source@1498.4]
  output [20:0] RW0_rdata, // @[:anonymous source@1499.4]
  input         RW0_en, // @[:anonymous source@1500.4]
  input         RW0_wmode, // @[:anonymous source@1501.4]
  input         RW0_wmask // @[:anonymous source@1502.4]
);
  reg [20:0] ram [0:63]; // @[:anonymous source@1504.4]
  reg [31:0] _RAND_0;
  wire [20:0] ram_RW_0_r_data; // @[:anonymous source@1504.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@1504.4]
  wire [20:0] ram_RW_0_w_data; // @[:anonymous source@1504.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@1504.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1504.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1504.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1504.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1516.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1504.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_data_arrays_0_0_ext( // @[:anonymous source@1519.2]
  input  [7:0]  RW0_addr, // @[:anonymous source@1520.4]
  input         RW0_clk, // @[:anonymous source@1521.4]
  input  [31:0] RW0_wdata, // @[:anonymous source@1522.4]
  output [31:0] RW0_rdata, // @[:anonymous source@1523.4]
  input         RW0_en, // @[:anonymous source@1524.4]
  input         RW0_wmode, // @[:anonymous source@1525.4]
  input         RW0_wmask // @[:anonymous source@1526.4]
);
  reg [31:0] ram [0:255]; // @[:anonymous source@1528.4]
  reg [31:0] _RAND_0;
  wire [31:0] ram_RW_0_r_data; // @[:anonymous source@1528.4]
  wire [7:0] ram_RW_0_r_addr; // @[:anonymous source@1528.4]
  wire [31:0] ram_RW_0_w_data; // @[:anonymous source@1528.4]
  wire [7:0] ram_RW_0_w_addr; // @[:anonymous source@1528.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1528.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1528.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1528.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1540.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1528.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_l2_tlb_ram_ext( // @[:anonymous source@1543.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1544.4]
  input         RW0_clk, // @[:anonymous source@1545.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@1546.4]
  output [43:0] RW0_rdata, // @[:anonymous source@1547.4]
  input         RW0_en, // @[:anonymous source@1548.4]
  input         RW0_wmode // @[:anonymous source@1549.4]
);
  reg [43:0] ram [0:1023]; // @[:anonymous source@1551.4]
  reg [63:0] _RAND_0;
  wire [43:0] ram_RW_0_r_data; // @[:anonymous source@1551.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@1551.4]
  wire [43:0] ram_RW_0_w_data; // @[:anonymous source@1551.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@1551.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1551.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1551.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1551.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1563.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[43:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1551.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
